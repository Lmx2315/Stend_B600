XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��
h%�b(y4I�Ϥ�м�2	�^l ��%j�g����-8��'��ѫ�Z�T�5�s�*/4��́U ~2�С���`M�gQ�6��
M�#�4S�~���:e�����k��bC��vm<����3��CL�����Iwzr��_��Q�鷤:����H�V�V�~���X�s;�H�Q=�~����T8������'��/�	S���S�O�����8�y^#��(�=�>7M����Tyi�%�a�‰9�|�x�G���%�[;y�?�{}��!�$������O��7[�)���]�o7�hu~���39�vYHwCR�<#�հ�=�N�ԛ���T'��&|��a�K�?�g��<�,kY؇�©P+��_��X�"��	� Գ����8J]F-�k�*�����u����P����DJK�c�x���Qˑ`��W�����dw~ �bwX����G�j�Q�?�m��z���&�����v.�u-�񜎖^s��;�}�Ҫ�Tڞ�����PY#f(F��ȗ����#u��ּ�PQ�0짽�m��K�1����� �?��k!Ct�|Y�+����"�C|<9|��K�����來��j[;8�h�J9yŬ9����r=	0����j��o��0%�-`�fEM�
aO�n��m��q�������'-ikuXsd���{��ć���ڜcn�ئ�B�х�&9�iXo4A����~�+@�IXԁ�XlxVHYEB    2864     8d0y�F�[��D"�]VL�h�"+B-���Y����[O��N���ʺdެD�+���*J��i�T�~QsQ�!ƪC��C��)��Mn�m�/�3V�o��6Eؔ��T>�S�]D�_��鰥�q�h� �dS����W������Ud�s�/����"�uΈ�MMR��
��*�_��z|�9���	6��L���M(ZT���.J<�ʾyko�@��O�r�lx�+������:�;;��߄SoK��B�MG��7��x�}��Y���0m�� ��H���]G�L���[�prp���"�&t�B�١`X�6�Ņ�NKY��x*J�#�Q-���Ý��E)����������-i�m����� ��A3%�l��M9�r��I�cS�s�d��T��;i�s/�Ҥ<M͂��7��(tV��tf���r*�>A����$�:�n���A���Ȱ�����q����) ~��Ho!ğ����i�$��l]���Fî�պ��a�%M�=�MY
6�U�T"U����c
s�;�^�Ru���I�D��0L�����è�B+���2}��eϝ;�PPE������)�u�K�N�GF�)�7I��P��Ai�jۃY�Y?􆦈�!ܒ����\2����<x�D��������t���g��8=YZ�`+\�䑑'����wV�ƚ�9n�0��L�ʑf�0�v�vp�e�^���*�.�^�#}7':��1V�֓���6[bU�S~F�����}�vd���]��7��F�Ke���{�-���]��u���p�����k.>}�s�Z��5�q~M�yW@[3��r2i�f?��A�o��������AȒN/��;�R�n�;X�^��\�����-����g:�B�������.>�Og�58��!�=S��,�,|��h`�X+xϻ�hV�p�j����$����y��/{|�OY� ���O3���:NY2�ІuA�ђ��Fݡ}53����"�d\�|u�	�Z#�,��Ұql�^�o~��x���s����1>��{)�ʶ�K!�x{�\&?C�6��hx���;h�Rx=|�y:X�W�A¶#ݥ!n�]��+R�I�3�B�{��5�k��,���A��/4j.1 �Kg�Gߪ}�Dlx�4���"�,XR��C���5PQƥ��L̫���ؑ`��a��\�/vk�2cX�6�N�N�%��dD��� �,�8��÷q�+0�ݪp�&TQB!۩u2/%���On\���n,p~f���Up���\�ew��It�����!�g3ޭX*t`�����3̦���t�WQ��@ȲB��28�+�]Æ�=�/}�ѱ�f��	}��?;��YVދJ+ۍĘFQ�7���F���o��uqü��_F �m�p����Ta`�����;�5+N3{aC�Y�5 �X�T/q(':֮����G���e��j����d����@���ؗ3�}7Ҟ�8�2d$��M�������0�f�9w���7)	#0N�A��#Lh ��^�N��"j�K{^�NBL~*:�"�ŧ��U��A��-oM���NJL��A=��d5gL����W�2]����z����sj���EZ�^����U�Ef�*.�د�E�GYR×��k�W@�m(W_Rfp2��0���A�Y�y����|��_���P�C˼��w�V���>������D��'����#RJ0FNfx-�;��]��r�$!N�����z�����F�\j��Z�>mH�)�JmAM#Z�w��}b|#�݀@ �4a�}�:Z��4�7�[-Tm��ވ�I�8Q��b��\�S{`�Oi*�q��^AA���� s���'�������vm8a&�J����36�pEU�0��ŭ<�<�z[�	��P�L� k���a%��G W*�˺R�K^JO�t!h��Y�ױV*` ��֥�ދ��1�᳘K�I�NB�L���tz�rM�V=Eu� =B	S�1NV1�Δ/���vlt���'W��C��A��àE�t��m/���8�
3�%Y�-�$��w����
L|�=��n�$�,ȍF��"8�r���T.w��E�x�	M��*�RR�O��s�޷�2���ϑO�:%�g��5���p��^WI�-hbB(x���0w��2+P����j� ?�'�g��a�a Dm�uB���]���ݵ~
��z��,�Gap�?꒓