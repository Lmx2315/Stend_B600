XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������̅8��@��^x�o��[n��)�9��ɀQ�����w]�H�c�vU]i'z*%��k��U��w
�e��>�Y�����Y�c]Fr+�9��~5M4
���e6Yc��$��ڬy�$�;c*�Ě^boIH���( �	�G�|�XV��qs�/ R��E���Ș�wh�����|v0��t��;Ak�Eɖ��=�4:+ƃ�����n�[�}VI��j�=�/�?��0��l�_��9��}�=V�!<ψ��4��d���=�E�G��1�.y4�T���p����o���ˋ�9�[_�0�/�K]�����d������T]�N�f���@��f6�D��Q�y�K��������U��T�v�6�+׀$�2�����O3w��4�h�ښ�a��&۳R�̗��cz $�q�eNi��5�q0�n���Ji�]��>:�x��K^�TI�Da1����x?G8��7�ո��klѥ�=Fc�C���]�d�-�I&�ލ�i�S��G�_7{p@\b�?����D��1���Q=.���t^�<-��[���\i�ݡ����'�`I ��v�F������M��Af~�A`<0��{m����$�_�?�<�[l��: �9�n�$����@1H�\9�R���W��b�����2�ۺ�fxO
ު�U]8��8�e}��=/����r�x�Ȳ��Y 	^�M"�D4z�ᛌD��hD3tI�䨬R3���sἼ]A[���_��7�G�yd>XlxVHYEB    1cf5     790����:�¤Qr�˝�j��˼[�IE�O|y��ʶ�#�z� 4`�#_ìaLk[�>`�S��B���������|�E���_�u�ȴOߝ�d���'�����1b��]1$�Ջ����'�Z�V��o�G=�}��-p����[�U��.�}M�� _UE��m>V�>�Q!�&����}8wp����/��B��,QXJ!=T��]��j0L���ǀ�]R]ԓ�� /��'��s��;$��H��8:�#�1({y�3Jq��#Ud��{8ٲ�̤�IdP���������H�p8;t����
''&6L ��T��P<I��j����mB�>���-�p;�<�Y����aV����I�!pz�ւ���
\�v��B���Ye 1�I�j�|~� �\L�Ⱦ̇Ug�ܜ����Q��48<a-\trm��Q��i�r�9�����$D��;!'?ɲr��W(7�����u�Gz����Z�2X�bͫO+�$b;�͕2��ӱG�Ci��\���~�D�\J;��g���|s�.h����65��ߣUL�F�B��s�,0�N�:�#(dr7�(�H�[[e7Ɖ8RʪB�s��0dJ�g���X�6�]�-5�P[J���$�mOЦ���˱���SV��Z���-(��or�*@�Gcn'%�L��y"�+�h���5fI/�BY�4���Z�R����!M�O��p�����7���!�����G����­��5������},�,��D��5�5��<�o� Z�蒵�tg�{�[~l�B�w�L��AS�&;�Ё�G��Gy�j���-���I�]�QZ�����Jr�t����STT�@jЎlѕ(k K
�|y���vM O�0Nͤn�l���f},~�b<cfq${r����'Aðh�_�z�� �f,D���Ln�s�����������`�m_�L��Zg'�ܨ��+Ժмq}R�g(9&�^���Q��͠��9%���,�#��Zahv�]I�.��^zD:�i�I�K����SGyѷ�O9o�=�r<�)���?M#��=���-�����Y���e�"����A�د�A|�'Y�`&Ό=�$�cmp<��l�����v�����F��ڂ�����1��!���Y�G��jU	z����V���=7�!�h�5C�v.@s�:�&�Z��+��mne8nW��p�P�M��3��C�4Z����(Ƴ��������Ȃ�C|��`����0��\��$�����	ͼ����W/ף��ѽ�+��^�a�_+m�%f�� �����s�C{VVK��k�����1	q��Nм�bH�m���ƭ)2Y(%�]
A �T�j�=�};Zr�����ؒ�Vy��_MD]nW�y����t(yV�~��S�����y�;�ތ����q<W�UyRn�����"���<TN'�����ZQ{�ߡ�TgA������e�2�@��?'��}tW�2�Q�n��E,2A"��c|ҟ2c����K"�y&7���O��.F-�o����S�UQ�]��@���T�|���H�8|���m�*mXƵ�U������d���Őc0��S'��j�������;nJ;�nG: (�$8�_�ݫ�8+�i�������o��i��+I*�&>s���o����r�X�ZҪ~7��q�j92e��|{�_��Zd�i8Q���4"�n��1P|e�@&�ݿ�+��$y��S|2u�Ѡ�8�D�g�'."ڞ�clDcI|7��Y��,\ڔR�m(�p�������Kh?F,���Ȓ�lnns妎�����7;)�[n� Fn]���/%ʼT�½����3`�p$�y�Y�+���r�Xn#>�W'莉V`�MsH��ଥ��@�M~��1�I�P4B��z��i�U=�