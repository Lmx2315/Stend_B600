XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��J�h�c���lOU�V)]�R;qZ��]ݫכ�E`����g3�jT��N8��f�r������QeY���']����)����'�r����2�������A���P�rL�%OA	���2�c�~�7�U��]~��G�ѹ�����=ϐ��p�368$.q<��:�+����� �3�h���{��<����j��Mo���M�x�Eo�6i���z5��3c" >E�U	Rł!�
�r�Yv���=P��@�4:�M�O�>D��f��AF����,Z^*�?���uP0�i\�H+m|�xa�3�O����Y�v��$�Qe���������p��x�<��xI"[��?(r{��1]'̖�w�de䠂-�?ѷ���$�S
�c��g�%�	n�>��_�1b�o��R�z��Ϲ�������H�|[?�r�a���.�]�م2���p�)���K!#p�K��p[��WSV�yCc���J�#�+��}���tC���ԧ���}�t�4�Z��$U�8���K����b���d�8�$�j�镧��޵�>�c� �L�� ͏I����S��{�-�|	�B��ܷ�S�Ѧ�|A
�N�i����3�$rT:+?m}Y�R�����:���߈薃Ul.
�`�F��:�Y��h3֩>�ڞ?&����r4D6���tgաH"�TX�Xo#R�䖱�TN�� �Ln�F$EE�߉5�4�>�.�������)��^f6m7)w��d�=���'XlxVHYEB    2863     8d0T�z1c���w�gy¸jM����
����О�hR`G),�Ko��,c�����_ê��wT�K:��`Nm��szs�����lb��ŏ�N�n'�����o0˼"���t�m��Ȋ��ʚ՟hF�Z"-�@~��z�}����� 6ka����E�M|�)�?�O�V�P:A�������Bvs��K`�s�b���t����	�� �Ӹ�Yb��r��9,L��A��)�G����/6��1Ð��H�;
��5��`�_߭#�rf����hV�]Jo��B\��.2�N� x}F�%Yf\�a�����<L�/���?��TL��rG�A&�1٠�ΰL�� �h�\tͭݎt�BW)��^�Q���.qu2��n��wm� R��C0��)���]��H':���B�2�TE�xp�y�9�'��3����nb�`�T���\��7�5�b��m*}��5����#��M��K�		1����N��p+rI����t�~v�g��v+w\���V.�������Sy)��8�+`�0�������	ynB�!� ��fwJR5l�\�(eS"Dj�x���q}B�M��'��;Mڼ�Ŋa��!�]� N~��j���kC���hW��蛨��2Y�U1��g�;o�N�{]��v��cޜ�lI��	*�oD��0�Q#�B9E�L���HV!�~���/?�[I ��-��@A��?����_�kȱ=0���3I�q��Zi�K�����ƨ

��Ui�!���}� $}R7ι���SmY��#<��&)A2���l��(��k�|���?�խj��X�c����=t+h�u~�>hGS0�� ?́���5r�ܵ��M��E�)II�v��������F��ۡ��Wȴ]_����c�Zbn�L�	���g�`:o���f���$�L����/c�;�z�r�!j�mTo�OI�ݪq��k�/P��j����}�~r�$T�f�3^`�8���e>�$|�o��O�m���$��0,�i�oh��`c .��M9�$M�a���g�#��ζCRmC��k��@NØ8�[��肻�G(Y �
'�`��U�o�LZ
d��дYg>�l�rY���:{ƒ��=aΔ������=�ф�Q�䝵�3�(Q0;����kg��A���]�~�f^���XS�@� �q*o�ը���bbF.�� �Q�/6���4�#����إ�>wͩ�/L�:-ް,���>
�!+�2Ғba��73�&��I`���&���?�=	;�*,�����?B���2�w)�p�&�=�2�W���rH��,X�[u���5�i������0kD�,/�Ȏ��VT4��j�v��w�E�&;�b�|/��u��?/�2d�Sa6f����U��il7��%�|�G12si\�N �X'/�����/�?��(��B{�������X�j�{+���>�,�����5�N��\VV�$g~F���U%���PJ5�NFc̒�A�ˊ@f��7���<;yk2$;�=�o�(��cQ�ml�6��P��J�&��fd^)�5;���� �$G`41,S�@YC���/��%�E9��(+ʹ� (�L��m�������X��X�#����x�w�K)��-�Z��	i� �lEr�^̪��pV�C���ңé��7m`�HTߥ̤�fS!9�ὪY�����Z/�y���u�҇�v�(ԑll�N/o�P�u��&��z��0���gw%N�Y�%;L�)��HQ[X�A��.F�E�o��S�I6���dK��Ğ�3%Q'dN6��?vm)�%���u��S͜.o2H~��E�7�څ¶qf�/�^��d)��<_^H�_R��E����d;R�������'��u����;��C5M���4$����� 9w�45M�$�LƏk�bim(��ޭ9�d3�>0]K�>o�@{�)�J�
^�{��tҦ�J��t˽���k�I}m823\ּ��z���,��@�MO�v�RsAԊQ�q�����&��[sd�b$ã��iD?�?F��FEP�=8�m0�V{��o 8�1#�˻L�`���Ca�T5����тm��gVZ�l)���pŊ0-b���#�z,��{�rN*��w,X�;�=N��,C�J�s�#���'@Bl��h���m���ZG�vn���f���>������=R,��gD�0��}��;� k���`�𕳃�م�X�:�