XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����Q��6�w�%�柎=�xj"1f�&�2���.z�5v�0�oz2J��,n�ϗPQ<?V����҄�~ܢz/�b�����h�Q��/��E�<8�6<Y� vH#��y2�f��j�Ф_����)Q �8�Y"�+`�׌�̃:�y4@AJ.�?�{�.����f?�P�P-B�"f0nP�ݥ	S��ʌϱV�QK��/_~�Kl
[y=��:���1�����x��m�[��fWce��訮2�_@�˺$i;�I����^�w6m� n��ޖ(�Eσ
m��Fv	v�	+�!ex,Ƈ)zl^����~	4}�'�(� ���q��`����r�����E�\��0x�,�>F�7������a�ti��b�g�I�OʋJ�dD��9$���Qph�0�b\��)��J�}Ў�|��}EJ0�3�_?�F��[~�.M�>7W��󍤳p����(����nd�e�=��^��!a���k�o�p�a\E�s�.��	L���V�eH�p�ǉ�D3� �I�x27Q}��M���~|87�h��q��{�2N�*;�$u)��^��7���Ȝ��[9=Zf�k��(&�Ut ����`9�
�� �_��1� ⅋�ӡ�M�Yzv��׳is'�ѺX�r�lPx�FzA�쒛�SN`$m�:o7�/i�2M���Gն��Y�;;MiU�9��,�a���O�����{/�̕;����V7�p�b�ʹДh����^B��}�~H$�U�T&jcO%�o���XlxVHYEB    3541     ca0g2�:� �C;���	Bz��▘&��O$I��29�D]3�>&�ww��)�+=_��P�O��}
���h7�[M�od�#��s FK���y|n�P'�0c���aߺ�5-<���7X�"m���3vg���<�4���]Y��s��H�A�X?".5�p���U\��o������8{�q<~H�<P�&�f�V�7$}F�7gÝm�JF�{����j�b�0'����Ʌb!�>���`A��I�߃5���D���i�+`m~l�썽+y}�7�:�fe�,�$Hf��I��r��' 
�-�O���k����9<�搗Q�$x82S�,�w��bu�l��@�$�IX]�Hr��2�Y���;j���l]ލ 0k��E�O�.�O�r��[♳�̆> �9��ZH��f49N�iij�Zw����z;�U��Ow�ƍ��r��џ4�2�KM�M�=�xh+����O���~$�l~-��5��g�q8��c�3/�
W���[78��#��$#T����"&�an���	�O��ȳe��nyEV�ƣ���xX�P�ɇ¨��ق�&36����t�l�]2�0B-��4m	M^}�g���]����AC�w2���._���p=z�)n�)ۙ*�W�H��F�C�()��.#󋓌�t�∄q�!^'����)��'��b���p;0�C�Cb���/�>�bѸ�!������.�H��� ��A
����v�_|�fq��3����Za���I����h��KZ�"8��<�:�7����1���ݕ�E� <�R1`�D�<8)j��������R��<F+a?]�6̞OĔD�{?Cw��sζ&����)�.�j�7&��}^�+c�̷zď�8����4��&��+>1�l��N9�3�D��P潈�v�������)~������������^�!���H
T���S���B�;�f��`=չ����5U�w%��FP3w�C����I������+�un�@��5�����֠�S�$�둧��[S�W��B�b��%|�	�H%�A�u��}*'{�7�~�i��Ԃ�E0��p��	��̮����Iׅχ�(�#���W�]8�wG���JBB��$��+6��Y�}�F�|�Ol��ݨ>���}�fF�0��QM\eu�)O�}�P&�E���oA�dNl�EW�2	U���&&�<�'�wtْ�(j/X�=�sy� %����?���|����h�>�P�wI�<�NvؽN����ְ���-��q������=�wT���Xy4�����v~��BR����i��Wf� M�M���,���X5��X����gq���S+=Z��$��Q����2�Sw�K�����/{�Jx�!�܂wu���8&`�sOa������	D.|���`
�3���f� ��H�@���ѭ�<�j�2�<�a��t�����B�&�5~��B��{�y2�BJ�)�u�K��u!����Hv����is����RZ�G��ǰ���G���ºa���Q�X�4-Cl�c�g�ɸ���c��/���U�����+1k�E�)4˺�e�9�I*,N���d[��!YϚ�vyݒ���N' ��6F��EDd�@�{�oCƠ��~[����A�0q��lq�/`��!Q���?��V���E1d������J�jAG:2~0P��ӂ��v�J"��YV	,M&QG�>Q����>��_�v$I�c(���$�f�,	HRyn�� �]��u+�� �.j�ne�ʿ���.r�ԃX[d(3xZ� ���U�����̗Z�܊�kE+L��#��cT;��c�EE,�;F�&�T�D`�w{�r2t?�4�	�46/<}���s+��N���{�ŔP@6��X�9�>�Q=m�6��,ɏ��fs���n̨�v%�G���_��L2zOz]�zWE�����9�9e����4��̱ �h`,���Ix��d��x����C3�G��Zq��}Ѣ�vN��L�F5�8M��2���Fcs�����|c��u׃%�4Ft*K<"�1��%s}��Ԅ�S�N$��o�O�T�|��|�Z��>l�_���#K�#���ߠ̺o7�q׫�PZBز6Q\�hN�}6B�0T�>V6��ũ�A�i�D��X.1	�e'�P^�P��m�Gb�(Y�C��C[�2@�6H8�v�VȮ`�$[I^_>E��Cnwҫ�4�|�t��G�"��ȜZ�Ą �(N?��Ȉ�-�F�f
넩�`K�&o���²�I��y�m�|�=�������@��f�`��I�����*鿁L�778+"�;�z>Yf�%�=F1I:{�9���R�y��S�Z)#1֔oN��/-Gr�\��4�C{F�S�3���� F�� �E�/,gE�Yϰ��O��-/���4�d���bͳ���O�]��]L�?�Cl����P�Wyk�Wř���AA>KF60*�V�	V���p���B�
'(�Z�6^2�V���@�l���~s�J`�Z�􌙭����[��P2��P�w��w�/}��+�0Cnij=�j,NSqM8�k'T*a�ZZ��m�(K�ܓjJ�<{Z��ɪpB�p�Y#�H	k���E�5���Kq�������G���-���ā��
��$ɪ�S�W���B��+��y�7�hz`��>��z콭'%�?�+T�K8ap^�PY�ɓ̒�W ^�A�EC70��*��%;Tz;��@9j� �j���V�e[�&�7��\�'Aad	��>SR���h��2�瀖ܰ�,�Xr?�g�p�����[����ߞ��TH� }�ϱ�'�N����'C?QP�3r�m����gP�ˡ���}�mr�0������xy*�D�3HlѰ
Z�G��63j_��|�3GeJ)b����}�OZ���ݮ�w�!�7�U�2a'4+��ڈh���r�W�0�dA��6z�xځ�(�,m�8���%��w����4J��W���I:Ф�)�E�s��=��C����ҩD���8�F]Br�Fd��dN������)^x�����l�ˤ^Eu"����?��t�|a��Ea��Kہ�R e"	�j����tB������
�:�7λPd=�Wi�t���Ծ��k	���C־t��8|��9�iݏ�1A�e��@�9*櫩2
S�����0:����