XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��^U��g~-�����iA�k�_r򴩍��v�<GJ�*�'��R8�f4�`Om�̏�}پ����[����͌�� �߅�ӿ��"�Ҍ#lJ���$�p��! m����Þ��,+J���!;�Mif���\r�f,>��� z�{g>Gd~L�!�_,d�I�'��M5���D�-�*h��FQ���ztW�;sH	S�hu=?v�.�%���a�9�Ri}�&N^���d��-��-��i�e�4!��=є�Uߛ�:'�Y��qZ����F����5���e-��/�#p��a1��J��JV��o���߲��g*DfJY9)�5�v����9�to7A��N	�a$��a��.MB-���h�'#ip���p�<����q�U�~��l~�o�:����my�r=����_��x7?�qg�q����Ej���-qs�ʋ_� L�˪�}"J+����y-j������,+��W��t3ߦ� x��O�a��U?����I�1���2���z&�k{E�	�Z���ɲ���^q
�����	��閣�ݨ#){Z��t��O,�uƢ��E��K�FA��w3���6���ee�&�R_�v�t!<�� ��� �c�?@w��\�G����Q;u�~ �c�U��:�.L+��+��m�pli�i, Ł�W �M3��[�^�1�qo�EˑZ^ L���O���s1���I�����Q@Д(X��"o1�M3k��V�ɀ�ug�w�L�����2_0J��;|�XlxVHYEB     b08     3c0Y��U��*L�����W�)��#,�=�/��N<'�yTP4��}�7��@.��u���.��,چ�`�w�Ÿz)0P~�/��8^�w�(Q�ᑞ��7)6Y��P�Ǽ<��b�[7�����9�D::3#t-���1��l�Y�b�h
Pŕt]���Y����]��NHn�69���������$ߡO�	'��}�|�Z4���.�Q�܏Fئ�l5c�ʶO	�W=}b5��~B�R}YSGR��(�p2C6���N����e���!&�S]�I�V,��{���		�aɯ���Q��ZN��c�xS���7q��I�9F�um���й����B�4*+��cM�A?��d���e��T�LS�Κ��������w��Bi�~h!��)q�:&z'�ũ�4�/�����ywϡ��*�q�!��-�kN��/����%�(CQ$���#�}$���߲�M0S'�
��6�ޯ��@y$0�̊� ��m��֕�������ڱi��\�]U0P�mJ�� ɥ��2������b2�#Z6�y��3���iT��e$7��I�%�҇x��_�_)+�����a$D���n��{����I�w�o%ˡƌv0�NK,.���.0��`k��<�0dK9�c����F�I�|��*��J.�x�s�'�}a?��ka '�yX���`��67����K�䴞�9ТL�;|WD��*8�H22��a��C�xe�Ǚ�'F͑{��s��lF����n�*۬����,n� C�����a�V"q�Q ���׿���e�\� �K��g�@{�bWV�`fpj|<���o��=��:+m�=<�%d+U��(��h*\	9"�f�3/�qeT�y��k��'�gMu��Ba���ڤ��PxM��ff��0U�I�<(#��C#�������q�e3�	;��R�s�HU���)۩