XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��eG�.�����EXkZ�8�nC�&�U�\Uv��7�fDu�z�ڱ
�`� ;���
9�Da�0t��~Sq��l�am��ZwJ�9���t��Rf��=�VĴ�sr*�\\z���lvn�3?�7b\K�xk�j�4�����ɀ�xB(ϞɌ�zJ#�g���>D�G.C_4%�}�z�G��N#����u�	�Vl�V]H�ߍmB(vo��$�7�g<&kkb�b���IW�3&�k#ፓ�[�)�|���f�S��R���(������*�;�B�2����oQ\cZל-�J���U����>�}	�Xd�K����ru�F�p��Ի:����V�5����� ,X�� $�C��w\j���Fx��͙箌ɫ܀MY]&���0Y�'�!��o"�fR����)��c��C��ebv��x�W6�9(JR#�N@��w
ls�ub�[����)#l���B��lF^l$�0�}4`_�q�ό�!ܑ��e��䘡-�"�;=_GK�c�8��^���645F�[�qT-���7\���U eX� �&�K9���@a�|)�o26/���gh�ViԀ���J{���O�E��6=�Ѡ��)�a�ztG� �ެ�]o�ʳ�q�!ʅB:���2X\&pXmW�V-����@?�_*�^����<>
�\�}��ߨѵ<©&��
TZ�p��S�lDNc6 R�j.��Ë�ȥ��b�7IP���|�0����G׸�çF�o�!Qb��>������EN�XlxVHYEB    690c     b10��:x��O��\K��@�&nB�_l"�q�qN`?�tQT1V�&t��^�>��_RD�p֞�t\���-P�چ�t�#
��$P~,�ɤQ,�ZKy�^[��IA�w_V��^P�C�:'��I�U�jD����񀻻B�\�������M���XJ⻭$���:Y��"B��io��P�yE��<խ�ʟ�G�����9t4�2ߨ��K�eE��p�:�s�E�bQ�]�:j���C|K�J���������>'��1+�{K7�E��x.Ѩ=�tkQP�S���'���.|^�Aq����QΪ���.ǳ�4/0o�!
d���=���P��Ϊ�H�.���+TC\P�J��������V�D��䁥z�K��$eͼ헂���p�Ӱ��mrZ���d�g�1J��W!}-��V����$8��K��dA;�~��V��llY�{��}>���J�F-zf��COT��:ߦc�󂢸Dp#��#��v���ݗ �s4;��KVs�@,��tdrz���IM'�	\iT�k���\)��Z�m�A��L�'��K�u'��q�ub��?��/&*:��>�ҝ�c
�H����h��BL]&�����9�\w6<S��3�B���q��GG�y$ƣM���3��u�wr�%8:}$YOgP� K	����(z1󼰊P5��%f+)��l����J~� ���l�*ia�F�U�2J�������{h\��ɉ!��]>-� �z�ǎ`�tuC��oh��H;4Q�6p�~��{a�A�&T7b )��^�T$i'�8������n9�>�:�:
�u�v���$�h}��)j�ꄉ��_A��F2(�5 �p�S%��I�o�)�j%��p75��]%��s-P��d�B��Q�%�cGu���ja�P���(I�liio�])��>�5H|0I�o�G��g@�`bB-0�4�xs�?+�!��},D
T���j#�#a7�����gf	=;�Q��8�n[����,x��X/�_uT��1�*D�o��Y*���dsHs� e��,�jo}�I��t�1�zR�/���C��;�#��/c%��q���N A�	fJ��C&ф�q��׌�c�N;ț�Fi��a�@oV�"�\,�!*�k�%dZ�T��00�b�2�P�"�V�յ|��m8,e�n3��?��0o�&Y� 1���f�3U8��h䵠Gl�u�(�	�#��]7�b� W�[�|p~��S�1�u���{����s�Y�����x��;q�B,�Uo#��S�8G�1�L�4_M�W�P΀��F�8�.���}��J�
���2^"#4�H���T��(��5	{R��������C��$��d��~��6�$�צ��?i	9�M�;�%���
�M���1O��$��&��u�6�p� {�h����a��p3�UT��207� ������Z5Q��F{�	���'ux���-����*��6�J
�x��;u�.�d�J'L�Y0�p3��8��Q�-D��*;�̂d�NSz��(���;�G��P]ew�*02�1�C��r
{碊�V��"�q��o�W}��㍩����1Ҹ�c7v7f���\بXȟ��d�j���6�����B��vه�
�M��a_�N���_/���t��?g�f\�z:�Z�Q+ /6��( � �I���qq�m��L����TG:���R
�o�ս�ј?��鳞�^��V�Ɣ55R�����q��Ϊ��yD��{1VO��AFو�P�ɞ��i<�vQ�(��e�<fۯ�n��@�{�@��G*2�ͩ��L�Ͻ��y_���� O$M8�5R��[���
0��{"̦}�^���+�p������ʮez��dW�����Ȇ	�gݱ���p|���D�ˏ�[:>BL�n �[��z�PsZx���Ѱ�YN|�TΈ�+�D[��W7��2�y�D%V"M &=��^��ͮ�O+f����rD�#��O�iI�g��Rٔ7�r��k�!���D�����R��x`���˅3[y�p�6��)��Ls遦�*WY���=�2�bT:A�Ȋ*�GJ����b�">(���p��]��k#bc���t��Y��ć\v9��� r�1It՚�����Kn|�f��u쇦�M�Q�M�};3��Ɓa������K,1��]��˩@��IDk�LCAH���
���Mj�G������O��}j$X�����4��1��7G�]G�^���w[?7�����V��f؋�1�܃�!�?�a>��c�����a�%���	P�kMH�l~͸��'Ā�ڞ����IL�3J�	L��W��/�����%�:�R�c����R��Lyj� �[̓���`�՘��B����*��D���N�0H7q��V!��������NS��NKc��	�>��5�D_RPe}��(�.:ě���,��/|n� �L\6�y*W/��;Q�ꪁ�4���pQ]��gsFT"fްf'O��*'��qs+Z	�\�0�B���.x�h� zu=K	o��{�m�U�G-Wi��NJǩ�W�Ŵ^�!>�l}�_rd���=q�(�����{6pq��K���i⪗��PX��i2����a|<Hӽ��q���Un�Aj�|J�����ǯ�f�f]~*д%l������c��o�R<O}�,"/����ރa���r��֜{����$�V�s?��n��Ŧ�R����0�$X�-DI��a�)|�0��p7�' ���9I�QS���;s�&r��Yo	٤vG�Y��5���[�}ow