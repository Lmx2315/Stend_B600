XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��:J��V�	ҥ��`�ڡ4�<Ƒ;��+� ��W<pI�q���O�W��;��+ lra�J��D�`�x����M�Y�:w�N����tx�����[R��o2
�a��0)������	��6��Cm�to�3�&��X?l �N�DMN<
܎5R��^m����<��`>啞 �@!�aHn�Q���d�fWU��m�3c�II �m0����>�n�1(��`������+@�Ja�Ь����-ˤ11�uQ��F�%Q
|N���5
`�v�����j���y���ͬ�����[�8L{����̬¹�����"���k��Ş�Y��w�7nǫ\BF�]ޡ\��A��ѵw֩I����!��[J�:�xqӀ��ɯX�D#�?ݥ)ֈJ�4����+ѯ�l�&�
�dץ y��@͞���Ɋ7��0(���,|z���k!�c}�]�,B�.f��]��
Y�+1���TN6��|����u/'�O:��s*¤�4M�p�d�m0�@A��֊�{��]Ǝ�KQ_Rzte�u��YMW�6���m��g���J2�I*[����v�� &
����8�\�)\���i9�f:0XF��W�Et���ܮl2��}kH�;����Qe�ρ'���d�kLgDshՕ�jW�x+���8���a����S��<>��+�R���q��L��
�P _���ёK���ZA�r�/C����݇ڎ�e�����b�ǝD��EzZA�t��hR��7/w<XlxVHYEB     935     3e0����dL_5r�|�&밍�*�Z ���D$,�6fؑ��pt�� }��3H�}�m.�:�ѡ8�zkv6��xeI��[���ͳ!�ܧ��4�53?gc�����\9�o��Sdz�V2��C��t�t:�wtr�׌g�9���[[�����Ap]��CK<dv����țe����xM�����^y��lD�\M�N�_�?�JC
��ux2ָ4��ߍ�&Z6���S�G-/�C�M�K'��k
�G�텚�j-�ԶSN�g������6x]!�W}�e"��ٸo#�s�r3|���F�P��v�B�#��F��	Ƚ-�d�;̈�>�n�����/qng�in���]q���ؤf"r�"�C�.rm=��ANd�<uvDWt�%@�f	k�r�� ���Ą�~ּBE/�L�*��QH �Ϻ(!��	��_Ֆ5�
��-kƞ��Zk�E�w����h>1pWV)ٕur��[�&�y��o+���N��sꙌ	*����He	����"y�L>�y�pϢi>m�>*�3j����Ԓ�u�;���w�n�s����.��1D���_���PA��?\�:Mi���h�>���,��Yemak�#��hQ�5K.��1D)�uJ� <���� ��rĊ	��V����s�E��]v���x�̡�O���Q�|�VIxeM#��kT�>�j]c]���v����7���c��0���2�����,丢��6J�����v�%)n�ė���Po�n&b3���i���fb�*�����v�g.
�*ReҺTa,a��<;���Y� .t�
�,� x�|1�n J��ij[�9`]��{�0?g��_��i�!��=�f�E��3�
4/����w��W������Fw��Y�5����zK$���n�'{��{�lIs�'��?���E8��@Dp_.zL@+��豩���W��jc���'
2FlѫKG\�R�m�w��	�Ш��Z��<ӏ�n��.�