XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����;K���IVs��w���ȳ�y67��Lv%*������oV�o+v��/K5�S����1�"��垵y��""�f:
=�e�ƙ^��>q�E>=�E�>2�F�d��{y���P�쳪�n��%0-K��i�p,��KJ�vg� @D!��Ca6$R:�>�G��{��o�a������%���X����x�(M'X�lN�L���������#ݚ���t�$:K�+���%Ij}a�>�ܳ���7Ap��au�qߌ24�21����C�#X;�3֧^.��?t��A�]X���@�MB������Ũ�����P�#N�-I�R}��h�}����Tw��Q͘.<*&�?��7���Z����𷒸�fj��/Q����B���;W*U�-���Fo��m@ǐO�0|���b�0�H��+�2k-$�|�u�v�&�_t��?EH��1m�Λ'.�	�_��-��%��*���@���#����J~�Q�+J��Ԅ V���k�y�`�����O!"(��6Uh̠�YLA�����Me���h����elZ2D�\4ϜL�}���
�2a���=v�]4}�V�y��̫�_�=�-�/�y�n�Ͷ獼_$� f	��5hÀ�en�qw�Ӝ{@`f8���L�o��'�3�闬W�K1�|G����WN�2h쪏�+�;Q���).��o'B�?�{�(�k�-L�?n�>�O{/df���P����1�1��tŌMO����INN(7+���o�w�e�q�.��`������XlxVHYEB    3a19     d40����>��w#0rX;�&���S{���ބn2p��&���)�)CF{�A(�ԅs�s<~����ϱ�z�G{�\9�_����b��P�B9��ܘ CZ�.
�L)�'��%�Dא�A����#v�K>@A�1�g&I2�-	
��|_>��l|��S�5�=��&f:����9�!D�z4�zr:� ��N��� �&��R{->�y�!F�@�U$�2��`��fTxNjw":���������כ�_�ă�j2�.Bpw�̠f�R�H�N�^a0O|��x�
yi��YW��Dh��d�*���h�/:�?���&l���@��~���5m���	��������Ȓ[�*gS���B��Fy͜��o龕ڎ�v�.P.s��y����IU����6�ڄȿݺ�\�lw�c*��7�f@=�0����n��a(#�W`�`C�Wg8�f����@�2�Ŧ������!�Dq�D����v�\`w�۟�w�~�����;��� /{��~�6��#����on�=�{�f��]D���'��3�]gn��r�/�N��I��T�[��~UA����$Ws���[��2���.��A�^�C��Y��I���4B��ŷ`�K�@�s�Z}9�r�5��<C�7��UG,���d{=�
:�ct6w[������lb�7�����-��_��]����)�w�NB���[6w\͘��e�y."�#M��-��eT��l|��;��<I��N"�jl��^<���3���s��V�uD�v=]����8��i��jj�e�⅝,�����Ѱ��d���υ�.�Uf\�a��ї�Ť�(֤�ޞ5uh���Bz���n4��������:��~։H�Ҭ��i�#��6����A̚�r��C�{����\S����J������FE�g�G�ƽ�3	,,c]�o���T�Lm�ǿ$hT��1j2�ܦ�JM�J�Ec�PBo;��x�b�s��o_�B������1q�53Ŗ�.W6��1K#�l�-��KZ4�\�F��*Nct�uA�-�ᜇ3�a�r���1��ӓ��0��?�<��شjuy�۵X($q�mf�����HN&�� �a�t�Im���$�[��H�_(^|5�al%���c�f��383�	b�H�gX�h�H�:����`^���_Ybc�u����?uw�-�D� ���#��qg40�����1�S�ܚ�XU>0dX�-�U+|Pv<0K�b�?�����+?o�	kc��̵99,�<����[|����,p5U`���,'�!���f���a����#���짒��ށJ�P���C�b�7m��|�~V���&*����|�>K��g�ìSRVm#P������D����_T�Iw��~P�luO�`�+~#DU7K�Ʃl{sS�(��r���������K���ʇ|�t�S �sa�F�i��:H�.*RQ9�~�e�s�\7��_H��]����&40���H�v�1~<����6-J�����W�+P�H���h�-@���2�� "9�t�O9lX;y�gkD��y?S=�fT_�jsoA��Y�n,c�Ez3��n.��O�Y���N���o�K���EpG�]���u��B]�WS?r��W����H�y���%0�KjN�Pȃh.S�:��m��is���a��۬�֌W�_Q���hyyC�E���:�iod߲@+�]!o]GP!,�k��|�������ɻ6�+G����G�NwYea�8�.���A���̍Lk�v����"�M�ϕ�-mH��A`��H)����BN�߲1����e��2�X�ȥ5�0_\bk�1�	�~��(�� �#�-��/�%5J�dY������8���C�u������V�� {�tΛ���"
�C�N��v	$��݈'s_4?_�i"����+����θ@�ަJ�e�*_짮���P�����+����SĦ˙��螑(rkDXH��պG5�%3u[�bտy8"��|�Rz��)秌2P�urNa�ۢ��'Q8�;|S���(�_�`!��3�ś��6d���W�gy�LI�&Z��$�+o7/��k�A8�w���ip��A�kP�lЗ"8���+O�\���Ɵ{�y�PV�x��V���l�&���y�'�~���t$|��󈩅��_�8�aQ���N���n�U���r�Q�h;V��5u��ʩ���zn��z�^�
�\�=�>"fx�,�$0��$��s��&�_$��J�lk���]I��oc����˛)�u���;�!��{hh���O��L����	}JX�O�U�Y�%Nf�T������ץ-��
Q�H�����8��w���.���h�Gj�.�S@[�)%�Y�h�t�@g���,+Pit�w��;�U)����}yb�wh+���\1�����k�Ь:�=�ͫi�]���jy��fB:�_��ߚt_I{2�h���H�.2�9%�4��[	�Ø�뛕�|���W�'<��,d3��J�j���ؑ��΢ӘKj��M�k����WA�eTq�`�F��=H�ռ�*d�����0�'��B�[�d�^�l��QgT�Z(�� ��M�I�T�U#��sA�o.�$�q.��ծ�f��3�S
)�(k],����&�b�40���O��2*�Yl�u�;!@��I��;D5�
<FC������C��~w��HS���{9B�4b��?�ؔ*�Eu۲�
�o�jkᘭ��7��7֏���Yg`�A�o(ve|}�?=��[�L��7�F!�5E�~��^h���N�>�ü��0eWN��,�{���~k�� 4$��$3^GO��ץhV�F��T���-fW>��&YOQY�&�J�]Aӵ���Z�i��8���,�_f�3O-��?@�g��PP8�r�]au4x�N~g_�'Xf��n][�2]�#��W�i��P��~�����ʪ�fʎjeXL=P��I��x�E����	�Y��{��Oѽ������k��pOW1e�,�ݶ��É���w+��UXZ�ВB�{�Z)�����<T#M��x���Gxk��J3Ȣ�g	0� ��-ȵ�;�����qAA�l���c�Q��&�`�Hz4B2#�u�o�m����Ȭ����ɂ��������l��S,�I�*=x�oa�N�}�6�~h�C�R������������yyN����nኵ�ݳ�x�{���[W�]�2�b��>@P��E��r5�$kʗ�DK�Mg�w�/��Cb�PF�]��������i��n�i[������po�)�b�ͷMTz�5[D�`S��O^���9��&M�S�䐪�i\�j��E�Oh��[.T�