XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Y�g
�V�Q��dԆ%X�"\�_����0��K��X�"7��.Vx{>c�6t+�w�ԑMjT��q.�|{钆��'�k���Jh'?;|IZ��tf��[(��4��,��lm3��l��_�e�z�vLq	�)\�m�.w��?x�l���ܠ��R����f�y7����J�\T0�c�oi�;��S��NdC:c>�w�97yIV�ő�(‧?=������a����}�#�-�r(���ȗ�O�'�V��	U�7)�u��L˩�Vt͒�V0d��:���ke���4��jR��g�OI-���X�+����*,9O�9��Bp��,��@Zo8�#}O��+?3��")�R	ωp[D�g���:t//Kk}O1���G/t�z�]�Ӊ(m��t��.��L����x3�Er	fM�/S�)AQ�ZC�� J��r���g!`@�C\��Ze:?�*�>)�'F^<c/��G���f�#���V>�Ɂ���qjo�E��Ȟ� ���_#8bBZ��C���GPs�)P�88C}�y��&�gP�����]^��v�<��5/��G�d �2Y���N��)?|�y ��F�x��W\X&���Q.�R�):�ٽ]k蘞�9�����[��%����Rn�6=Ħ���� i̼e1�׆�݄:�]�<5Rm ��D�7�Q\G��%�c��W�8f�a����é�^F���rŗT�	Pz�?�	��P�+��Y���ɿ	T�CT%�,"@�5:�n�b�^�V��9E'�XlxVHYEB    1620     6e0����6�����^u��g��O��rx �^H_�2��W^�Q�����j&�e� 1nVfq�2E�s�sH&��#~i��A߅�/D���D������F���+͑yנ���������J)O���~�
���g�.�te1�}؉�z�7S����ɳl�TG�I�Z1�̺,Gz���O`� P��T����D��؁8*��5�݇�q��pz`Y>C-y�c�բ��A8���.x��_�O�`�ӼÜ&�t�l��i���6�yk��jp������ѯһ}_��m��J�l�Kl��v~6C�8�T9�~�qG�H��'C��zo�\�-����<��md��x��C^\�M�w�#�Ǖ�,��0���:����%���S��)\y)E��0t̶T��a���duf��s�s
�ㄫ�u�H6��dCN��ā��g�9�!0[ӡụ�Ǵ"�|u��QFՓ���=�{8����*�gw���)s=2�?I>yr��E�����"��4��u���|"p�������-xe�S�C,�,:?t��Vy���0��V.��S��m��{ǐ�{K��2�pc?N������|�q��R�G}}�wn%���~��>�IȨR��������2@QmA�ӹ���uQQ�q��$����icí�Fl��Ju{�MW���ָ�M��]�o���*���qÁ�
�������썆��$�٥�z�s�h�F�D;�sڊ��7��:M؈(�;C���i����d�-���
���Fէo��@�r橨���
����gr���@�n��J�dR	��2]�g�G�qO�y���TSA�(L/��vJv���ȓY��'z�H�wH/��xi1�yz� G�x����"���աp ��F�V1s���f���i�̱���؟$�U!��I.}3�w�Wo�6Q-x 3�*~�E;F����=�t�	`~�2b�qǠ��PC�!w�$���[ú}�6����јkO~��*�e|�W�>��<�n
�c	���C
<4���y����t�4 ��h���<]g��N͈�s�?{.��Ĕ(\g��{�]��,����d =%���=��p���>��-4Y�SfmfH<Nnɴ�V"����5��(jI��0�$#�`�� u�߾g����[�4�I[���g>F\[�1BN�nO�g��� �v�	�rkV:�}�e�p�֏QIM�ܮ^@ګSt��Q�E���������;�$voa�zN�7Xv�Z\wi���h�Y����2T�C�~���δ&M�`&ІM\I�y�M�c#��-O�n��Zޒ�>i���!H�R�xE����o�K�Ki��uX#.�t'"��.��S�
���ItI��Sy4Jq5�L�Y�Ye>���
�(�VZB�	.#�$�U�Y"�@"�� o�E,�Zw�[eg��l[�[&��]\R�-�Hz�^���2�-ƶ���F�p�0�� yվ���ɫ���qU�6fWJR��^��K��7f�Jo���?�M-�Ti��(8��Bh0�qd_�MM'3���&�p^�@Aǡ�l�/	7��<�Y4\��!1����u���r&�(=�Y3��l ��������HwMx���օ^�s0/m�����/m�;̾6�J��bb��}���o�N���LR�y�	�V>Bv�1F�ep��k�T���(�zȻ:)8cwy�D� H�x�<$�]���m\���Z�L�a&lE�(/l�