XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��;��VHꢋ��2���.�^�G�X�X��E'�4���v�)��]KP���(����d�����2��K�w���oT��CF��$�_��J�˔��k��.���J���ȡ{aR��G;�A���[GF�d��g�����!$�_B�Q�>y�-��sG}&�`�$��w���_�f���c,~u� �8�%����a�!�1F����,&m�@���l����P���	8=u*��H�b��Y�kѶ�8[:o�3n�\��p]Xe�ݐR��Y���_���9�����[^��P�Ci��r��u�/?ut{��P�Fg�X�ڄ�|Ǘ�V2U=�5�GY�s����<��Gd���;��$B�#�λ�]���j�"��6��Ў����	���9�/m�������o:T�Q��L�*7���'|��&r)5�^�a~#�RKt>N/�
����qu�5�}x�>�a��T�%6�>�6RD,�Ƀ��Y.����Uc�[��W�͸�@**h���Rt�L�O�<�Ka�*j�~#m2��[u��>�Q/��0���<��'Z�T��
r])�1
@߭E*�."Hh;hJ�ޙ���,���"a�S_���� ixݑ7�?ֈY���/J::�<�=п��r[��e����xoT�El=E�m�C�7>�4:��OЎC��1�$k��Zx���2.-�"���7)xH�N��U�/u5�J�B*N�-^k+�7�2i��u��%Y��t�j}���+�G���%\��.3���@HG��XlxVHYEB    1cf8     790��0�VU�[+�V�(���������G�FvM���v��{�od�>�d(�3KgR2�,4U�_:T�[�
<�s�ZzO;��·�	܈�q9�vf�b��X��*�)���IyJ���|!L�l�Б�7.�/�Ε7P�vt�u  |�a����>����������y���*�^>�_C���p����%�.�)��j��w�!9M���l�+z�A/ew�K��B9(|�?n����H�f�仦�&��#��Z���'�����藸I#	�\.��r�s�#k`!�
�c��+6Иę`�v&��WA=�On~C�_�O�ɸ1b�#|�㿿-Ǝ����e��re�����0�NA�+i5�Q��s����\"��^E��e`�v��1��gꮮ^?�1�;����1��(X@���~G�%m�9$�K!�z{D[J#$lP����$ɒ{��k�����U��J�n�M�����o ���5�.ÉX(�DE�z8���+ ��U2t.�=)	����E �>��
�O�ȡ>vMRX7�JcѶ?����q�rH�FH����t��;��V���y ��b'�XJ�	 :?o�y�Ȱ����\�	޻%ꀕ#����ӫ�W�)���� =�H�+��:�6T��h)�/�VR��2G�$zAӑ]�&C��fb��l� �	�V9B�����t? �����ɮ����U�����D\)o�7n��I��qTcX���?��A�/��o��7�כ6��� @�[c���:��ml�w�K�=�gz�\��Q�c�:N(�Y��cY߰+����z�`S7�lܛ��2%8�={�'����TWr����b���
{)vvZ�rA�3En{&f�5!B���П^0c#o	x��l~[ T��f�ӊD�N����S�=��,/\��~�c������t����G��%sb�)���c�>LNT�0E�����j����PEM]����H��rG^�Y����V
��gM�V�'.��r�i9~���SV_ڰ�M�{�6َ;z�=p���~�j����5hG�i(������ӹ_�uW�I�������{�J�%�
3T��o�_�ۅ�!�J�ᒋ�Tt}��,CCh%�VR܆D��XW��b��[�1�+eŇ�:�sf���>��lr.:�R�1N����Mf�v����uD�0�d^d�|�;t�c��D�&w�ɛ�/��aټH�{�D�2~̻V�	���݉.�|�Y� %+3Y��U���"gptȱ�NT����y������|ʝ�o{u3�p+k��?��ݰ$s�5~�f��٤Y� ����h_ì�=<JZ	#%;����jnvQ���w1I������d�>�,���i�h����PV�3��d�>~(�?Ú�uW�n�K��P�����{uc�	p$���<���gY�'d��d����*< ��� ���a�t�9�}��C�;�z�[���M?�n�񻞦�/�`�6D�L2%�X20�aq�^�/R�E�-/�^�s���)��wn�l��(p<l}e$U6#���r��O�KPxz2Bj��b�3)��B�l٧�p�� t��3.�YH$5����>��$뤫s�2=ϟoh>��O��¯3����K�я��M��]e�S	�]�^wU���FdMnh[�����7 ���K�u��y�r�������옵��u�y��F����a�b٪xHhY�rF؃��)ѯY��ߊƚ�>B½:����xL���d0�*i�$�t{�:M)<�X�d�# ^ħ�e���;���Nd	�7b</��1��"����!D+��8��gZ��m_G����uUe9�s߄�,O�n����[l]�DG������L8�q o��X2愇��w�E#G$\��YJemw ��F