XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��_���x̓A�'���pL����nE����ܔ�S0�	܈��!��N<��:���$:3��i�'M����O�|�И��"�h�QSw���1��f�F`x��7yIf�!�Š�?J7X՚G2����)y�9PT��w�am0^����\q�i�r�'���$�t����eCR�f�t�E���+7x��"+�I�D	[y
iû�� �ϋVb�]�`����UYqh����R�(��v�6�_)U��7�]�l���0Yx
�f�6��gn�-y��>�yk�]~]��K��3�6��M��B��Iٛ�1�l
p D�I���iE-�]m�%Y(9E�'0~}��֣��R�.)}�mߛo���]�+g��MFYs�xZes����vBc�H�!������8�#2���_��	����*9��-����&nY˚j��>��$*�SG�3�AQDc�Z��Qm`�B�pVePq�W3�(%hX��V^$aԒ� z����ʿ$v�F0��X,ٯR��-��^.y�l[��Q���sg&{v�����4�����a����Ʊ'��2�_�� 1oI�Mp.V����AU:ƃ���
�"�~L�B5�ZY�i*�	����.�4U>��C��6ma; �S�a�/TP��Rh�_�h�Z���5��ׄ��Ka�8[|VK�J6/�`��rO�B�,3��S��LƷ�W�
�L4m�C%�5��~IJ��pW���2KĻ���À�����O�*6��u,厝_��e=���XlxVHYEB    1cf5     790r���>�j�=�k�x��,נ���K�:���8�2��3֖��������n�wט���-���ߥd_-�/�[�z��d�ը��m9rg���@.;�ШׯR�Ɵ��_�-�"�ghd�}3&.e/_��y���@RQ,��|j���SOT��A@5�i�3�*Z�:��_%���qm��~�x6���6F�<��xV��9�P{�IY[<����d�O�~[���#�P�|�ݾ0
��y'Q�_S
+R]q�v��B���o�Ѽ^m1ِ�5E'oR+�˄qA"-�O�?ۙM��;`j!d릏�.�Rx n�!���qv�`�<�QX�/s�#�]i@�"w� ��P��Z��<��k� =ie�iU�1*~� �r6�E��x}<��F��(,ʉi'VA��x0�����M�Ǳ�s/9AF[�=6�Ugcv��\�PbYPr���8<��"�K��Ư(j����1h��VG;=F쨍�ae��Χ��ܬ&%�zIS��KQ;���b�ao�pg��K ��SO~�i�~t���)*;8'�ɼ�d-/�GX&�6C�q쳾������N�U��W����}� �.<��r%���M�2��� ��98���ʐ�R�%]�F;����&�g>3ED�e5"Ox&�y����f^��e8��ӥ�i�����gb#q/����OW2�v�I��g2��%�j��Ġ4q	�M��yN)�q���X�kK��j�7兛�@����F랦x�\	�������0�z�<Ys~S�p1��� Y֜�2�f8�� ���c�j��k��WȄn�D��v�K��O��+s����M.��;��g"]O���Ӗ�L�����TtDs�?;S���	���w5_
ZÌ|�m��ؽ��N�!e�`��Gi�ז���Q�B0ԛ�t�B���FG��h[�N�W���52�� Zf��;��o$��8Rˋ�&��������\èf���bpw����ZpQ��kqi��b��\GVXiFqضK�%*���#S��ɝ�a��� ʎ%[��.����f�P�˪'m!�����+�C;]�©�ty�V�n�����.�Q<H����ɝ��Cd��4�NֺR�M��b�p�V*���O��#���N�O,Fn�"��AnЊC��Җ�N�ұ�N:�N@�n̍ZO�*�y���3��dl͌ł���aT]��ք�E�ȃ#��rU�P�	<'�OA��N�q���-�Ví��%4����ֽ�0��_ZE~j��4������}o�/ ��%���49��٣��A��;+�+��%MEq�DD��g�¼|���i�Wz�}7�\BK߈�E����e&��T(7q+ẩo�?��HF�`�o��\&�j9��R�s�h3ٖؐ]�঱e�¡ |Č^5W�.hr8��������Z���ܑ�!rJI�� ��26[rG�H��_��;&�=�ڈ��Y]���ڄ�l�L)AT����W�#�m(,�QR��d��L�����EbRt����C+�eK�v��ތP��|��з5�Y��Q�̏��{0Ġ�
���t���"��4dn�����:BO�HG�s9lv��.Ҡ�PV�]L��+O�Ig_E����ڼ~���e9c�WރuŸRe��.r�Ր��s,h�	����S_�d5���9�R��)�O���b���\�?��~%���k���m� v��F�)���^b���O?
l#yV��~M�[�2���QjU=���쏓�8����f�kC��6����L��I�k����'��*�,��Kw{�=���#^������LQ��IM�"����%k�������G`q-c�d9�1�*l-m� �&��Ł�ͪ��ǡ�:��c�b9�ֳי��m�S3I �Ƚ���q_5�