XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����(�Aۻ�R�N���?Bk��ݲ��:H��	M��Z:��u1�@��Dͤˤ�����t�����{���!�^	P�@yN'#�8~�)�4��'�\��;�Й����ba]t�(���n'bw>����!{x�(z�G���t^�Γ�Kܗ�NE�S�sO1E����K��T�@YY�\��	�QX/��'aWK ���?�8E��8�r-�Y v�
��:ɽ��U��?z���������/PT�k� �_9��M�Bcym���$éiy�Pfa�U@^;���vďrL+\���2�+�P4�����U2 ���+w�X�Ɵً���PG\(j>d��`�	��G�ҟƲ֭W?JK�X��i��y�^4��.�|� �z�;�Ԁ����`�g�K㪽K`}pqڟ�v��V�`�2��'K�����j�ce��{,�⟑���F
�����"� �VM�VQ������4�vOjK4g�p�*��3[�L��O�_�\Z���#FQG���	`j�_?�1��͞������Ep�so�Fs����L��x�18�U�U�d_c����ub�������������$�eaS�kr������0@d��n�&��V��Q�{9J�9���3L�[]�lq�@i�i���������=
�z7^���܎�r���ь�5"����^TQ޴���2�LDj��K$��H|
��FR�+�WԷ�^6�!��'_F������ {d�I��C����iBOɡ�n���f=���+I�mAsK����qXlxVHYEB    d88b    1610� �%�H̜9�Z���k9m|���=�J����cYP�P���8��zb���$��I�!����dp��Y*�Guwr���-��/n� '#����#��IP��s�*����},�n[���!�C}��#�4��1�Q�"ՠY5�c���ޫ���5e?��{�^	���!�m?��L��0�����H4���L[=��E��w��Q���[�ٱΡg2n��2�B�a�1�!T��?���zڒtR
�3���ͦ��\'O��m�TK��1E=5ۡ�K�ۀ�
��a��YI��ܷo�³��J�����?x]�gf�Ա�8*�8`e�f�y�	�.>p�Vv��`ęj���p	i�-���|��t��aӫ��c��?5��p��޸��'rH˘Uk��ҷ�_�s-��M�L�%����e`��^�tL�m����ۆ�g��1�/t��V����Xp$`����$��, J�g��	�r�N2z���4��3�^�ՋD/{,��ދc�4���#��Z��
An�w1N��D���0��x�Ae���Md�ne_H�x���&�@��G��P���/�(����Vx%�<0�� \���}��C�D50`hE.+�(� ���j>\�ɤ}�����@�8�|��4����G Ml��� ��mNa�a`�@���79���_��I4��/�#e��3�&�ɯ��l<�΁*`zy�)q� :�d��d�9]�?Џ;wv��+�(��Fů���[�3�T�^�;�`*��ى�#_ r�a[(&$�_̙HS��c��С�2	�l�QL����MY�#{�<����<�,(&�>�����Y�;0Ҿw�D�� v+C&���E��.��.�l�Ny�>����vžr�&a �V�Wp�o�ш��R�;J8��a��?�CBY��CΚ��-�Z��-9Ɔ\)L�S�R�9B���v+낶'
b����t����G���Z�K���c��i��Ԫ�M�پ6��� d���v?�������8���C�$�p�S�����,1�;���f�&+a 7��`W��q`z����g[���t{�Z�����+#���ܜx[��hVi��(<7嚸+/� �yżLt�Q峽�#;/��L��S�[��y/���b�$'0o��Y������GE��H��O�}�\��WH��# L��|WO(�b�x����L(�j��dg��U�$���3���<6k�=M)�=�
�����Ks*݁\-|ވ8Sq�󡴦|l1��ԗ�6KA���@XY�w~��B��V�L��h�nv�3�i|R4�����W!�g����+,Ju>ƍB�h�o�pb�V`�$wV0����� [w���9���]İ*��z��ҿ �&{�Ԝ�M�w�/����I8��v�������)��n�2��3vC�qQPg}£�x(}�ʝ�?eYD��*B���M�[�	��_��*�uUݔZAqV��|wgP��ˈ�)Zb��G[�yn�M���3`[p�������%a �\�6)��U�RXm�D��j��0[�*�Z���Bۙ-M�+�����MX���!�z� ^E�� ��>���L������=ؘNz�Y8$#�w����[�Q�@z:)~:
[q��9c�x�P����{�c������Pd���*�v�S����U�C��5{�r7�-�˲��tù�#��;�
������W�.Q�];���!i3����9��']��?��V����d�����6��R�-���LN��≘�v�Փ�	«s�q;,<�h&�H���Zk�����7~���tC��?�<=fn.�~��>��b�	�ku�d����*������2���\=�
&�;��݂���+P$*��?��&R{�(wF]����$���Cz��PO*#Ϟ�+<�	:�<!�!�� �B�ݱ[����*�6uW�FŦs!$L_�T���P�Gk�5���Uu���f����6�3���7��;�0��Tw����=�@]��f�]���E��e�b,�m�I�&��u�o����v��y�=M��
R����TX��I���8�g�Tِe�H�l���c�+`�+(��'.�i&�4L~�+)�E�fEO�Q���Jr���<>h 3S���#�ώ�̓$��D�cU�Nۃ!:O��W!mAԫ�N�%3����wfWK$��Moh��J����9g�
Ɣz��g7�DT��v�p&��|��i�5)6��v�&ib���$.�6t��Rf��pM�!e�=%Z��ʼP��`W���^-�����MҎ��\�"�n�����*Z��ˠn�9�<�J��{����v�����)�7��s�����)'��3XNU��r��k2"s�f��Rie��v���i�{,$�]&�
Z'&�E�B��k�^�ґ�<r��f��Z���G��W�Ѯc �*¶9��̓�H����1��<1,����F�}o{�r����k�`o(�?�r�L҈P"�,�'[���~� Ŋ�T<�c�qa[:��@[{�կ����<����"
�)l֖�J�9���T�뗼!���V� H�"Y��ԕ6�=�����R�`�R9Z��dj�,���2$7����>쬩�BA�QC�D�,V/�Ƹ]�Hf/�CYP�	u6�Q�G�x��Rd!�nW�PN,Fsqe��i %�v���/u\M��8�:e��A����c�Xһci�SR����Qs��aygRe���B����z�hk�����_p��W�3����<��z�<����e���ɣqM�tN�~v�ٴlˮ��:;���5��E�®��A�p`�!l%�fH��H��>��G��T!��)�i@Q� ���%�bΝ̱I�/�U�Ϝe�C���o�MZƶ�#��< �F��?������&l��|	*��*Qk�7�j��";tUW�C�P�eh�ҹ�ķn���+���9_�Mκ�c��� �׃0*ʘ�Al>#»�yFz{��^Ȥ��`k��<Ɵ�գ�t�+�� t���W��&_@�췵��S� {�����ȴ�|e�Y|CO�H�ʷ}�k��Ƌ�W���^�^�ͱC&��v��e���0q�u��p����#��_]{Z���vT��X���*�����b��1����|{��/��>p���r�`jh�x���Ib����&��,��B��1����O&{P-�>\�1�k��4�,|�8L�XGc3!p�Vߴ[�Ҽ?\�$��s����bj�l~c��T����MP/����g���$�V�Oo���h�-W"'�k�@vR���9ѭ�N�_L�;rzr^FX����]����L5|��v� �S�Z����$�rӯZ�*���$�RLM�~�
�������Esa�?�ie��W��='-�1pF�|I}��4��前�e��R�o���l'�7�;�ؽ:�؉T5�.���.�(K�6���dn�����k(#GWJ�!�B��;�s�.<yI0U�`䡂RL�W��T q�d��*ANG���h�v�C�j����U��z�yy8z��"D�7WN�.�	0A�*�p^4��gF�\��f��4[���=Ã��xn�UO���m��L��5n����ޗJ]nQ�{����߳�!B���Xl��P=��a�u�[�/Xs3C�J��ҥ$S�ѕ��d��#�����<���ۺ�M�Ӓ?3�����?�w2i7s��x�� "^~��ˑs�0�rs�:RA�|_��dǠ����_1;�VΪ����p/7���y�&�&�8����]Y��7ua�|B�Sa��Kř.~k64DugykLRNfq�Z0��J5��Zx�2���� ~�k�=ྕ�B��PJ]����0ʜ�r'Qj�A���V�.��\A�JWi�k3���"��~Dw��K����T��זq�����N0To��������:J��E��Ecpo�b2�d�F��J��}��8��l�\�Ih�Q)�~�R�E���AC�1\z��&��7��/��b�rM�L�n��jŁd�x���d|�s #y>�Q�O����Ŝ-��w��M���ne���Y�n��Qq���g�Mx��U���dt<� ��������l��|��b�{{��J}����gּ%a�����&�Q�ch����̭�>8�b�Np,2b}���<�l�i�M��sb��4���[@���x�V����r���6oVY���GJ��L�F�2H؀�g$��vj9�q Ά%_eD�u�W'�Sw]��)�녿��W�^3�I�U6���}�2K!�O�t��"K� n���ޭ����"1\n<�sF|�ps��Li+:���+#L�.��:N��L'����kcs���x:$vq�w�
�rI�_Z�2����c"y_d,�a^���I�Q�[��Ҏ���jW��XVPk�����t�, �,�̇��q��9_P���W;�|d�J �:Jc���]�hl� �~�c���h^�=֓�'�X�7S��Y�Y�9�2Hnc<���IT��£��c>�
�Z�g��v5�'ݯRBJ�%zE��aC
�L� #FP��݄���b�.�tr�2����L��ں:�Q%��UD��]>�(�l��R.�$�ϻ�d6���o�=�Jgm���߀&� 9�����=1�@$��A�H)�{��?�~���4ڡ^��[ ����!u�9J��	~���*{��6���|^r����G��SS��h�5��2�S@��9�0���O��d3��ط��~�`��Bk@Wu�񸶱�5q%�ѤJ�0���s|�&�Hu@.ά�T�x�u`�a�<��>�	|��fn����h�Q���ݞQ�@�N��:ieSA�8����,�����k4�����j�dG��B��R�?�Y�'��v(���LV�y���$'[7"��؆�}~�P�~�{�� �W��s�Tz=��w�	!�abB���G�S%�	�E����N�hoe�\��a#a��M����$[ڨ�h�mbʞ��+ɤbη{��ʪ�yBէ��{��~�Խ�a^]�XG'�i��&.�Tӕ~������S�����m��6T��(t�-^���+���W���.����1)Y��,R>�d5� ۳s{�Q�ۛuH7=M#1��)>�y�|fcrV)���͐a ��C��ty遫�O��jR���JG�2#l�X���L�,{D�.=����r �8�s~L��Z;G%�C5$����2��?����n{�f'�v [�=5�&�,s�!��j)	Q-�T�v�ç���(��'I"8�V6w��Lc3#�J�#����v��>->�A�ϑu�	�s�%���O�5p��TK���L���&�w.p���I��:ƚ�FU2nS�[���n\���`t�vy�R�P�������GA챃}����,B6�aJvp�H���$�8��a;t�v���A��~���cO�HG!�v�M�r��]7?I=�%����GS����5�����ϻ�b�j3���� �2�js����(�V�
���k]��'X�_�7�1T<�#+����5��8a �wA K��MR���Ɵj