XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��#��->d��b��I ���W�M)��]QX/J��$h)J�,���UC��<���;t_R�	���|b���y.�kV]?������]��Z@��t��8.(tie��#�,�| Y�i���;�����YK�Y�a��h����_�b��@h��@Ő@�{9�6�z�n�c�w����Y����u�@�kȉB�q��J,���d~���` �9�\*��\�ԘB�f���[�J�/�\����y����L�߯>�Gk�	�[����{�; RvC.C��4���~#�1z�Rg��s٠r��������gi.�Us�eK-�Z6��O�1	���}��f�'F$4w���%y�%Ǩ����6�=�~���(��?k�p�8��-�x�v�8:>V��\Mm�E��$`���Yҿ��N�U�F,���;��)��<)�����,Cz�3D�})���ˑ���������nޠ�����GK--���ӧ���ޯ�\�٣���s���f��*� Aq�Dj�f������ QZ�wz����Z���0�]���s��C�Aj^(wv�}=���r�|y�o�S���j�������=��>��#�����Dz������P�6�|��f��2x;�pmj-]�D¯��g�$�~5��ْ	\���J�sjP�=+BN���Yϡ)	���1}\F�������H�G���G��3	�#l��K9{� p*ٗ�%Dy����`���,�'U���<������XlxVHYEB     b35     3d0��E[���آsv�,v3�.J��U�	3�6�:Y�ϸ@�윌><�����{�3�!�U�,�;�ab��cU��w��=�sǂ��[nK�_Y���C����B���[��H4�gff��fYf���+��]}��y�������\_*�����k��[K��l"�`�
5�|+d����nݖ�$w�d�"���A�!�����T�M�M2��!�$�O�uҮ�>�p�̫��~�)�?�'�4���WA�7�w��gӛid�K��f�8�B�Jଈد�����Sĸr�/cՒ�Y��E41�W�V&���3���]�×$0 ����у�?a�J���C���e8{ e�)�Z�� +�|gAo1I�!�7j��� ��8����	o�V\U�ie=Oy v��������G�ƅU��~}w�wo����Đ..��B������E�t���R>5;c�G��,XǓyx�z��f�A�f���^n�U*^�ǂ�=�w�f�,68u��4�I��^E�l{v!�J#��>;�@���D����?j	)�^�����^��
�&�,rom�\5�`�Xav��-�h�	D��>H���\=�v��K��e��5>{���i�I���tҺ��9'7�0w`sYv�4��ܶG�T���0*ڂ��BH,�e�(a�v��#�ћi�K9l�Um�[�#����SN�#_u���%��F�ʔ�����'ae����[딀O��Xm���`�Dސ4�+�I��]�p��-\���".`���ݤ
1/��wO����0[L�@�qޓ��'Z-��㸠P�W&r��r^�a�S���r���η�+/�N� |�OTjeՐ�ɶь1�E�f͎k"U�^
�>9S��*���=`�������Фl	)����r���-cN#O�\Zc��	ǁ"�w+���P��E�W�ЛOS���E'P*�ȡ8������/R�f��~�P�h֩��