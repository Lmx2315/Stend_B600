XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��� @�!�N~��AMϼ�}��1[��P h#^����Y���cdUl
!�wJ����}_�Z%����蔫"�4E�,�wβ�GM)��VGC��h4�ۻOM���p��1R�І��?���]��l
p��F��o�U�S�ɴE�c����Y�jhp;,�F;]���ճՂ���VC��2��#��^�D6~�H�s/'�j���[�ݳ�J�.3�e~
�(�����5C�����%f��ah��iH��#-HJD3u���d��mgSǩ�(ݽф��X�{�9���j�_�//l�m̍�)�}�:�ӫ�G��%?h|z�+S�@�J��-;��$����i������׫y�~�4��,��ntW#M��.}�/��9ى�E.����R�/󪷭�A�Фĥ+,�I�@L��ox-1����Au�:��[N6�l٠�<"�PH򲔤�m����I���Ŝ�	�ȷK�F1��E�\��m�R����8��E��YC]�)!��@�Oјz��.�XqL7MCe�*���~��]��c*PMa�U��W,�}�;"�-Mg)��8Ř,���]��Hb�5m-��>�Q�KY�!{�ob6�?�P D�k�j�u,f���>��p���DR[��N�vAW�zy[���=��yP0�agƒr��	ޫY���e7҈Ԟ^���6��b� Rx��ְ�
�J�B�D�7������A|�Sa�
��R���˳�bbqn�x;p�o^�.��<�s�O�lƝ�pCXlxVHYEB    1cf6     790���	�sQ
8ܮ��x��f��)Bp�B�!ͬem7�4�E�?2��Z&LY��3�[Ţ�7�S�<�D�d��1���1����τc���+ÿTT�(��ƞ.�ն�v�o�8�ɾ��O񠴀�:���������G>��K{ӥ6�#d��[}�B�U��
u~D�-������@�To�{��$K��0��O.�:� (I�5r`�35P�ҐB�N`-рҍ�åWP�D���P��v� .9����N�g�Om�(l�7�u�)��F�EL���lg���H}e�����@۳4�'gs9��T�y��Fe<j�MEuݢ@�:d�CzV�n/ly'�*-u\ڿ����ꐶ�ܖ`�/z��xb���/�G�5+����$	 ���8��7"nu.����
�%M[�
�ds#��몦J�'3Rl6���ܓ���?$��D�\s��H��#�8����=W��e<Z��?D��k���>�?7�景�W�4pTW;��}����2C[M�ч�"1F��c���k�O�e駾|�0��_���<iυN�
�?���ANt�k��'����rr+_W^8�5��0����d,��B���c�9���Ash�A�Ż�=f֏`�2���8�nI��d<�iu�4�	+G��1Qc�=*� ,zt������wB_����i�[7�*�\V�6�h5_#�,�7���ߧ��yb~+�'�8����֗5zlM�E�y�_kU;���� ��-��PQ�`�гԉu��	��VQʸ�K�2�ц��op�Ո�}0�5}H�lI�D�v+��#�q�R��h�q̓��R�
���,�� ��#�E�,/�6�]셿�ں�����T_s���K���FA��d��aB��b~����{�����o�17A������vTQ ���X�>R��zbA������/�.:�W� MO���kՊ~1r$%}��+��j�m{,r!�:�����y}?d�ݐ�$�.7���8]�z��yN�����4��(1s�Z�����y�▖)�+q���]?Ӿs��Hѻnq��J)��uU��W�ʶ~�ny4w���J��l���J�6t���.,��P���i��E��K��:��Mx�ǯ��$���\W��
�� &�k
x�c�A;j��4l�6�sT�6�ͽBWm�Q-�ٓZW��%�@~pH]i���b�|]�n_R`h�*R��,8��3&���3��]�u�h3�hϓ��M+GXV��Ў���7%��Dj���rG��n�^�~S���sA�|���-8N�ӄs�C�ݍ}���v�E�s|���n��:d3�����{(�H�K��BS��8��DV!��4i�\�s��$�\�o�����Y'vލ�f4_���i/����&l�Gu�GE2�̪���[�@@�u��̡�U+�2=X#<G �@�����E��t��xR�ݙ3�qUX�d:�}����B�=���w�T�Wk�v�I�]~���Q�w�t�ԝ�Ƴ��h7�Vr�!�2׋��%O��u�m8��0�NʌC�ޅ	R�*�y���r�=���k�;�E�k5΍te��� z����Ji��NGY�h�m��]$k�`�W�b9Z]�92%J�8�~��۞�,s���(:�Q5�%.���"�Xy������X�Hw?�9ћ3��(`�������6�lߒ��5A#�!��2b���~��,��et�.�w�牺K��5�i�=��=�z�W�f�+I:ؑMCE�n�.'D!!R8���Ϡ���J�H�uN�.|d��C�����[�*��_xНd���Fh��oAx8��8���$��EM�i�/�DҮ0����*ȵN$H��}�D�Wo}h�FR��_�k���9�VhD�Uׇ��V���N��D�aϹ�C���$���<T