XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����|�]�N��1?�݆�ܐ�Ig;'�=f���ʤ�s�H9�6��Y׊ϗ����s?�5�z��P���:OZ�՗0�����!��%������z#G�E����n�F%������0�|��9�;<���X��x�gR�x��w��î�m�ЬDz�!�m�����kؚ���ro�i��pU�_O�P.�}��^�0封�Z��(�j%gC��X[�˯�$w�D�v �U��
��Ď��~�o���!�U-i̪S�f�\K��<�#I�K8��ɉX��A�F���M�k�A�����= �9�ڹ�N*˩dy��e���u�Z�A�������s�vqP�ǞOz�:��!�`�R��>y�.���;�^o��yhq�u�?�~�DI���f�EK
<����l{2�(���{е�){�p�Y��z���=@)T�ķ��z,VtƝ�'� K���t�3(�́ࡾ���G ��|l&�9�=5ߪ+�ѭ��2~+j�i��m"�*��?o}��@u�],���$ӷc��#�/��װ���ZCsX���ӑ@aF��z";�"�@�������e(ӌ��o�����N��_ fJ։N�>ʰE �
.�w̚o��B)��3}�Z��s��p���G߃����1vMYZd߲%4��m��q��y� �TᾦNMR����2wM�U2���\�Ө:�K�	��s�ޜ��O�a�mŀB���.��������M_�s��r
I���r�`�P�ă!^�E�mh����k�O/��i�XlxVHYEB    1d52     7b0���nݡ+0��g��?�4���ռY�{`�I"�pt��eUu2�jX���]C��~1���ǒ=��@OJHF} =���K`��<�8��#�?:ST��1˞H���٦��ޥ�|��!F`.r֏z���n���y�[c�����'�y���?*��ה�t�I��{��M&����<k�T��n
�׋����s�������k��P�ڝF^���̧3����jXf�M���c
�	g����>T9�c%ECn$ө�ay��w�iTQ���ٗc.��Nx����͇9�kތB:�Q\�7SU�R�v�+�P �i�I��Y���]�}��7I��le�Ԧ�7 ���3�c�pLż��B��i?O���:8�]3���S���o'}Hf�6���/��'�|d�K<��jV*)6��-O,��7�Pd�#}y�ǙyrH�l]u�}p'�0��L�&W)���s�	#��bQ7i�v��}wG��J~¬뒈=k:�w�8�ثg�i��-`/��+�R}9^��l{��$��qZ!qN6�"t򾢁��D����s�*,��|WѪ�ڝ��d��th�����Av^F�g.��⇬1��W�vu�D�`�%a�`m�#��SV�m��0�$<+ )	Q�K��f�J9`t�Ȟ{�C=�_�G�@8L	<�K�*��t�9��!yV+T/����b�W��9�Oi7�)*����(giAA_����q���?�R��q"�L[���"j0��F�{8G�7��� �1������kwj��x����8r�`��$X�&QD�諂�"6,���R��CY8���]:�ǵ[�U�ҏ ���j7��-a�=�}N�_��%I`"Ch�C�@�Ĕ�+6e�����|K��a����y:�OW�ټ ux_a�RZ�p�~�P	*S-L�k�i��H�j4/���,\{}�|fF�����Ks���VEx�}Z|)�e�p�E�c�Z�w���0`�n?!�r=�%W#J�ǎ�.3���jh�Oʕ<�˅x�`Y,}g%��S����3�V*��v�H���K@��A��В��S<���h�q�xE���������A(L�
:N���XS�1K�z}�����~P+щ�p��-�sm�:�-�Zꛂ-!r�1�� K��|����{  9F8t�DLd,/f�N��$����v��U-�P��?�>=톰uE�>IZ�C����JZ�E0�=��� �!�A`$��o(L����;�_����L�R�ۓ����'���I"�Oʷ֜\9�L��1��r��:�n�S�ꍎ�5։�Z�x��@����&�7W`��$V4s4��}�p\P3ZC&a�i�]����y�W:��%�����o�K/��/��8L��1�����~�: Թ�C�مw�㹩DmSέ��RC'}��q�8�N� خ�b��9vf�bm�$��F�Mb�� l�N�<pi���&Kl3�a�TH���p͍;:�|$<�����}@s��!}?�&	�*����a|�K��Xc��m�C,�É���L���揞�����])��D��
�z@�X9�&|�$u��Z�`��+�	��FN�͐���)ɇ������^�����gr|��rdb���a/^�y���0��T�T�*�:�_g��+���y�9�3Q�8.���\�n��NOTP��јOֹsؠ<�U$���ȝ����<���2�s��݊O�s	lΚ��Kd�G?q�k�P����|o/�������?����
�a��]�%D\"�W {j���� jò����s!�n��K}�p�z~L�腑��@��i�ʠWo\��N��+32������SO��Aր��+Y��4�OC�K��@;Y������J<b
�bD�2v?����umwH~���v}�u�z=Q�e�YM�(2k_� �!�G