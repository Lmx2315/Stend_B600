XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���v���	�V�V��ªU���1 uS�)��9igPQ����Zx}J�3 4����%)9�hx�*����Q`���"��Ѫw0^
x���yHTra�: Hʊ���j����Ŝ0���	E'�\����T�^'w&�UK���ͻ}��iQ�`*�|� �C���|ccf�EuJ{O-��ݣ��'Q���~	O��S�PRx���a�H�7�RE��^tׯv7,���n�J>X�3�q�a��(�%�$����jS�C8@�)���F�TX��B͜	�kF�I݉mfOL�S ��#P�QF��f��WRޢ�l��ɘ|�"f2Z��ic'kFˢo�H�0��_��2��i����i8��|�V]�**ԉ����M��W�E���=ߍ�}[P�8�X";�tZ<��9kG�q������P��Xach��`�a�@%9�DĒ<G�X��D�ϔ�DřFb;L�X�G�Sdw��z
ٷ(�t��W9V�K�������s`pc�ϟI�<K���o.�X�@�H���Ժ���I������=ni��A�pP�5>WZ�94��f5�V��0��Z*A���Z�B�q)B�Z�-@q<䬨W�QZ��	m��eoE:�,�k&�&d�Q�(�.�>U���ǝ�lD S�j���C�O�/SGL�����������%D�Ok����H��;����c<�{��AZ���đ[�wn��o*#�rK�BE���S�o�(���	2�:���l���g��	������XlxVHYEB    5a4a     590�����B���7w1���j:�}%� �ȹ�'��%g�l�o�WLݿb���O��0��a�x>n�����w�]mûosm��w�~���D���pȔ���F�����68c��N�S�2��J/���sN_�X=���}){5k�Yù��&\ko~2��i���9�o�<�9��a
�ͬXE��S�p�j����٣��^,Q��=>.�m+�urЛ��/���:�fQ��p��et�x!�����negT������(�$-��8�jI�`E�
p������z^G����%�kd@A�^��"��]ov�] Sݐ��Im&':A7����,��qT;����W� ��"���yȨyC|��=^V+"��X8b:�����0ʱ�����]���{w����[�eĢ@Ŝ3x* ��+�e8k���D���sd��O��n+��%��E:�OLЧ� <�\�2��l�C���W7�'�2�iq��F�p8D�%�Z��d F�?.&��~3��f�4��DFT�L|z6�\u�n���0���D@a�(���":�m�;��p�s�PM�����b�@^X1V����V�MKψ%�X��C�d.F�6��O�&��,C�*���޲=�
�Sf*	h2���`Ya"�ۤ6�D_E&��}✭0|�CD����y�E#�di�QB߲DH���pV^86�A'+�����9x�5e][���f�'/����$(Q癧�)/:���������(��:L��ҁkpL�:|�7b����8(��Q��Ҟ�������e��vi���(���E>�{�"C��r�3�^q��BD�q�o^ (.��t����E�Z�Y-E��)�ٳ���9�������^[����T���s�as�|pl~AdwQ����`@��e ��ZM��V��u�5u��R�)/����6{J��y���x�����<�
�B!X�Io=���*&�n����S�.bj�{c�#�R̺8Y�jU7�y�G���
�;�	��N*��j���]�٤̑��E�s�b?�1����C	d˔qZe�V/�����L��s1*yz �
�������9�UգT)�n���F�����0��_��SZ��>�_�ּg����16 �	�c��O��M&�7])d7����R��Gb�XX���N��Ŵpj0~�@p;�n�g��
��ijZ^:[)�<�3ۯ4^Mq�oF�P���c�	��RQ�/dF���B	E�9c����_����2裫p�n\�z��h�])���t"q ��ƣ��[�&AF�2�5�g���e�� l�� �> q������r�=���/�����/�/��RROCkj�s�,�5�lǿv��t�<�8���̮)��ݑУAt9\/!�VC���V��`��.��F