XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��"���HI�BQxMs ��w��9�W�*z����D]�p}@���>EG���t��$Z��l| ��ԅ"BŗyȊ��y��,��OrH��SZ��@H����ۛ2?&0:d��r�~ ��@���!���v��qܖ<bw	��.t0k�cyX�|��L�}#&�aА������p�<�Ϳ���.vk�%D��+����]N�)�"V=�t�p��-YZW?���[��f쑝8�srA,8��!�G�-B��t��-�.�7vu��'ƐZ����_Y�����W�N�ז�^�ݠ�8p7ؽ�\��N��LcH����b�o
҆�ǿ���lT+MD� ˘Y�o�
�I�.q�G�yu�R��0}N�ST�jEֱ)��D�Q8g��J-�\��f�>j�F#Wy�C��>����X;5t3�V!VR����H�����.�T�j��\C���`�;��yAL8'���i���<Izй|�����,�����_m�br%f��-VjkW�v����9>sWS�d�l�-~�֦=E:���bVY%Rv#�ʓ�i��ɋ�v��S�X�b��
15�bMKǯT�:a�FtVA�"�n��`,&��FH�	S�RF���@���pY$��l5�pa�/a����`|y'��j�t���/b@X���Q�Y|�
1�\^4P�#^Ź9��l.d����7�s�t�M�#�Ac`�"���Y���Ś*RD���^�5��>�R���I׊92L�t��	w=,���+pT����{����4���HhXlxVHYEB    1cf7     790���f�6(�7t�a}M�����Q�<�Ĵ g'�cF��/�J�.oiǿm�|�b���mE��(Bsս�Q��}*|:���iE���Ӵ�G�+����?Lk��Q_�-ڳ�?/8n�;�Hn�1�e��t�8�;�꼸ǽ�5�h�j��5Xpj����>L�Ի�I"����_�jq a�^��e���G��L.����K�#i6c�gU�r�DP�`7U�����{��V��{����.�w�[%>���E���2_���2�xv'epˀ_mb�Z#�R�E�1ﬦ����Y��ؘ*|`@�ܸswM���Q�gr9�`�N>�Q�8�CV?p
����Q���Q�xMz���a+t,D'Է�����7���=���HF�}��Vf���G%�:����.�E�?<�uD��MpkҴ����*��Z�����}'��=K,�.Y;�OP�돷ov;bWWQs�6~S�1�fI�]��%�nߟy���h�(m����WC�� ���n�la�e���%9�u�������q@�QT�j�I 9o�4�|L�Ϧ�Tu�(��d7
@��+���&���P��A����®�W
R!�����	+�+�
�kW�M����5�z��I�5�	�v|7�vZ�{73���1�.g���Ka���*���P��L12��ų��6�z���b`^ ә\�7�f[+A�*ro���,+��AB���hӞd�{]����y�~��|��3:LY6v$d�O���*3˅<wܠ����\,�|���SŲ��ő� �|g������0П�>�t"�h��f�x#�4����ot����F�i�Dp\��sCX�ľ%�	;�w���@��HXAA��Ӷ���ݪx_�Z'���/P��;�O|��T����2v��=R��!����A>�^	[���XT�=��L�w83��9��Cc�Z�i0�G����P���1ʅ\���
���c-��Ecz.
�����#Q�����(���,�nУ@""�i�i0���W���Y��Me�~07��z�!��3~/P/]�[f5��d���_�F���R!l�ٝ�G�P<e��d���=��\�D��#J��L6=Xl\:O�hNU?x9�{ޖ��(4�c��Zm��Bȷ�1w�!*z�@�kB�S�t=2B�}q*���(}�>�0�\����^��TT�e-�^�?/��ǧ�>?F�xA��Y*����\a�gT�=�j��z���7�M�,_L۩�\	�C�Jh)�R^N!���
R�ٕvSX�
��/5�IS�p|�ݳ��I0���H�7�q ��$�]�=bG"����W��Q��c��J@����D�U�L�て���	ޤХ�h�9S���PH�?��,�����
YL[���fx�X��$1P�غkAk�(Q�>��^@<+����}���XaLi�ğ�Qh��G`7�)V�[���UR`���� g�"�r�u��ŏ�� '�Jx��7���n? �*k�^(\��XMqra����ڻY�uzj���ÈX�H��}NRH�AŢ.
	RW���q�nk&F��ߗuO}AKNߴ̖M$l����
���/�`�����_J�.&�PڹDq�c4�Hg?���<vu��ğv�ߍL��f.'o��H���屫���
u,�F4N�۩���H��C���",���H�}�nɁ^�D�����c��r݁\es$���t*>����xH{y�Q����z�Rr�=T,��V�@C��T�Y��ܾ�Lj��_��P�����9Q�=�X��ո���v3�[[®d��<͊�����sr;���c�_������꣟q\�֒HU3N��F��c,@he�Uc�a��{�z�=�)�-��1���[f�<�TL��iG��ں��˕�-�����`;�Y�����]�