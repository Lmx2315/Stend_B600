XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Z'�cvp�~�ý����3�.�&/yF�'Y�.Rf�L��d���̼f���h
b+�)�H��X���䁙���ג;�
�;�����$�0*�y��0WqA���􎗲�*�fEu��ȴ
��x�95�n.5G�]!l��.�b�w�M/��^����ɘ&�@���I�K�����XI���Y9���
Lv=q7)��{����$���ѷ��Ѷ���ѠC�H��<�9��NY�}��jȷ���Ǟ�^n�F��3�l��=��wK����D �ֹ��C���T.
F]�w�D|��K@#
QrRI,v���$�!�۬J/LX��^�8�:ta�3�x<qsQ��:��bn��sf�l|�!}�������4e��eE���"\рwy~G
��l�uH|�	���g�K�QgJ��F8���GZI㙼�F�w~Ԋb��Ԇ荈*�1�A�ݣ_U���c�
�N�;\B�:�2���1�m�^oؕ�6��ۜ��lõ��ҝ�N5�h9L��q�=��ڪQcB�z�A��P���W�3��F��HdBI7H�M
j7�戗Z�=T�s�{��b�!��g��c���̳ΜX�x/��fG��2 �?y�
W+����	�������q���{�u h�Z=ߚ��8"t�����_���G������������]V�c�DN��:Y7���f9yKK��	v��IX
�h�m�K��"Ť��cLE쓢���~߭n>���Z��R���j�hOăD�ͥ!XlxVHYEB    4e25     d70=1�t@�\���5����xŜD��ib�P�"h�Jg,ӭ�"gS+*i��A������$^=�k�/�of���a�f�z5��'�2~�)1����p��L?fK�`���!�s7�X���愞�L�9�BC���`����������ګQ؅���H��E�B {&�����6����D7�;+RƳu��CM�Ct�<�Ŋ�sF��etv'���9�B�^���*�L�Ϫ�������v�'��k���k��R����W��dQ=q�C}�SKJ�V�����l�=
<��L�f��z0X�ʺ�P~cG�4^�p>ԯ�� ,�=��Jp��~7e�WC��NvF ]�5H�����V���i+U�2�O~'4�����	1�<�٥3M�<v����?�0��1p3��J�<EM�6$���0��MX��%�E�Y#K44�D�R�T�)3
�z����T@a!aĖ�!G+J,�p܁�Jv+?"��Xh�%�<H�"23Rf9�<��u�q�u�-3�	KSF���M��s���À�D4��9%;������E=�͡N!R!�U��P��Ý��f5��'>�%�!�������4p��.��~�}|�u���4�D���
���sk���G��Dא:�sv�-}ޗmsK����.;�k�l�1��O7�dz��c��[�I-;J���ѕ`��&>8,|�g�7��&Q?D%*������LaqFh����M���2�#s����Fn��D�v�Y����X��Η�g����.͖r�y8|F���$=�z�b��;���Zo�U�R♔��ʅ7j�� �1V�zY�M�L���-�1Ĩ�<@c�dm�J'"
2�!���˳Zm��^0�@�L� ��J�T��=`��g
q�~�SG��'�
绁>ZfL�y�y�Z:��%f�py��
�F�XĬ���)Mj�����{��M#nM6��2���qg_X�$f�V�h��Q������۬���ҙr�+: �0/Y��Bپ�a�Ro˒P������8�Q�4�~���ER^Rۼ.C�G]���.�v���\@��H�r�Q��'���F���'5t�6��=(�n+�WR�h���w�{��v�y�Ԟd���=1r5-���%��4�� �6:r|a��k4{�qCG������l�G�"-�M7�i�c�
N\@��⨪�n�i�me�;���-&V-{��&=��K������oL�];��j�F���a&����a��\eTz�wS���e�?��@�yc����L�ո���6��F� �){�e��Ђ�1������6��C梅=!���%����� W��~�R��^�k��*a��z`�"������/��=��7�U
�����Lŀ6��l�Kt���xēgEئ���>9����t\,Xǣ���'�m퀁���NF������W�Oa�5�=5�/�I��fg7q�����>!���h<���Dtd��gN���LoJ�2�t�"�@���E��Exi`��K=締1'r(�^��O��`=k:ˢ��ލ#������~˻3h���d��z���9-:��R�YTr�c���.�#����8#85���f;%@�emm錣�zU2<�+s3����"�	����'�������,�{��1^7Yr)�'lض���FF�
X�����f�;�b ��:�`4B�~��2�/n��@4U�0r`�����j,<��"��e�����s}SC��OV��o�s��߅�$t���A�a~G�Ŋ�����"�1a1��o���m�>2��vE7�[ó�#���<L¦���Y����}ͳ�'�ͤ{��%W<���`�_�&+J������3<9�OC2�
t�Rt�P�<huV�� 7��&�h Vg�t�i����x�F�!�ɛl\.k��S�YN�ZױV�k�k6�8L�/�µ�$��p�`��H�\E�9;�/\�iQf�E�H�������o���l�=['N�&�Zd<��©-�R�@�祄�]���;����6���st�{���_O�5O�eA�F����h���jAN,��F��L����D��M	6b[���\�i�^5<d�%%��ް��ޠ�eF���L�D�Zr�_�8�|�S���������kd"JL�l��a���Vc9w�-B�%~��o5�T��^����]\�e�V%��f���9ud�w�����A���y�I���z-���d�b�Dm��O�eJ���r՞z��]����ʚ'5Ay�	�J�=Pa��@������Di����U��<Ą`� c�jg���*��ˁS�E�	�DL�ǃ������`�b2��k�m �\- ��T�z��|Q�v�[��d�����e��T��i��D���S�3�dNd�1p	f�����TwUu��`��ϸ���V�{>E�U�`{��lɰ1)ŋ[�M�"�-Cl�>CE�r��[�/�%tѮD�3e��< �;A��	sx�/pP@f�H^_>�9��-9���dmb�������jV;�th�z=�����Nb�W���P֧�c��V������o��c�=Fhr# � ����N�3�E����>zUG8`<�-��(��'X��,V+���({��*X����C��L�l�u�&��#@���ڻ�ċe@���������w���瞀<­�]��.��%�������S�ǰ
����*�U!�,q)�֑�s��"�����]�
�l_O�Ǥ��Q�;(6�<�z0��]�jZ�!8�q�)?leVz�ZOm�����ߒ��lD#�����z��[p|~�ڇ�~�22$Z��� �x���x!k@jpz�;�B�T�����U�}��8�����o�͈�ֆ�̈́뮓�w�̊�G6^�^��=S��0���B^_���Z�4&q�S�~nI��Į�~o���A�vW�e��C�&� %3���h�]>&:f�h��Ĥ�9x"W	���O�D�r�~٘�т�gY@����k���>q�������.<¹�q���J��O7�ء�r�EA]rR��=��1�H�9�"����+ę0���E� ��-2�=�j�3�^���ߙ&�z���_j����|�K_)$I��������!��G
�A�O�]SDS�Z� GM��e��"{1^�Z�C�������3����t�d���Tx=O$?4�tO��l�@O�5������x먏�6�>�9:-�qN���'d��5��_M71�w<ݸ�e�%8�9�7To��C�	e�ra�;���;V�)p�T��W����]�ꑘ��W4we��#��������'�����b��Sb���B|Ւ�q��XHyw�w��0?j���W��`����_�DGS���������rpDЅ��SA�S;1h�:�Lmz��&�