XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��H���e�A2
_��>��!�J����ˠ*|���;8X��vb&��ڍ�		�_f���U��w�I����5�fB��l�a��4邖{&vd��|�~��hL��%�4�I��&��P�-��b�y��Z��O��4 �b]q_|FƔF��xOD�sP̭�����Y,o-f?+x�����5��!�fb��$J�j��\u���1 hy�%a������#u��0?�#Z~������eҙ3�ܿI;{�d�$)��`LAJJ? � �еK���#���_��/^���N{⎡�s��U�4݈y��|e��@���4��;�6�~�\��xÕ`�˽W�T�{->��C���O��Y���=��$;�"QG��ݍk���d�/?�O	�{�K����M��[���hX򼻯�(dV&�d
��t k����a#�-!�	��P)lq$� 7d{�a�l"���p�
��6>�ݜ��/�s�K�i�!�P�%u%����$&R�Ыi�����5�(���ʕ���@���Ϙ���6�
j�Y��D֎����WmTrj�4�z�;ǟ��]�
��oHn�%C7,r#��$�Y�4 �F��ɐg����?L8���*����K�V��Ո	�~��T�(:4*(�0N%��N_��$�w��DS��V�g���ƥ�����)�y�����b	 }�uvW�Ĩtv�ȗ��`�����0Co�+ZS AɈ,��ݟ8��6l�� ,��Q���ps8��l�ɢW�Wz0cċQXlxVHYEB    10f5     490�+	Mr�˞ĕ�p*�3FmV�X�8cJ���%�Y(�ۑ�.;=;�I��#�;{�Dq�sJ�1<�V%�*]w���h�E����ؐ��.F�B�֐(�,�	��Giq�(",�s�n�&�4�3�y�}���5@�H��AW,��q����{���ۅ;�I/D��V�;�ݫ:=�6�p�n�Y'�q�� �;?�l&�D��{��w�����}��|Q��^�:z�9�I���Q�C�m$�tX)��>d�V��O�W�g�#���h7~����
�灻A5K���s�#�����ҟ�U�:8�A�i���gij	�rE�W.j�?�Je�?#�$Rn�b!�v�o�8��DՀ�0N�ي����D����Zs߯�Vw��v�w�ˁ��J��ۮZY	���t]w�ĲlI��8j��I�U
v�9�;�;/!(��c�`SU#�=�zI�P#ƲY�E���ثF�kJO���G� ��nj_�5Q���]�9��]W�\k<�����g��A�@b����{�K��0�<D�����hrhWv�z�4z�����Vd�� �@�d�?�j������e܋�t��ʐ� 5]�7G�	 y6<59MK��m��֗7ܝ�����{璧� ��hѰ;DL]��̳d� �_0'�4Z�e��NJ�����Y�3�?C� �D?P�!F^X�l>��e��6g�b��hQk܌_ĝ`���r���dy]`�J;)y�3�Y\~�4��(���k�A�n�/�J�=t{ ��6ԣ�~����M�*�y	'���̼l!����`S�0�K������)���l�{"ԁ\�p3J�>vQ��]G����T�Y��.!a�h��lK����<���+lh�`-���B��F� �N���#��$����h�f�zmԮ�1�����E�
{Z_��4֥�O�z-c�9�y�wEu��FUcEh�jy�Қ��XzZ���q�M�j���=o~Ci�(l� \��[K9BG�b�N5�E,*Oƀ��A��PD�5��v�����Z@ʘ������8�Ut�{Z��Sx�h�
�$��~JG����[�ۑ�J���wË޴ ��dEݺ�A_���|�BU��6f�Wr�����/λ��� �nj�;��2�8�5@�7�N��1h���� �6�V\��A