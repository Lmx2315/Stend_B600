XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���:F*����w�y��W���O<��R�E��b�W�ȼz�.��&x�|�D>��2nsJ��b�Qq�K$��w�<x��g?�*+:(�,N9�b�����SP#������v��%���D��ё�W�,�.HV]��>��QGW�Wh`6��?��WϺ"׺���{B�)�f���;�1�J���7��;Cl�$]?�fPrF�9؄�w��f�յ.���x&eOY.�Ed�5���V6��@��t"��SĦ3gg(F�/#O	���=�����=$.�
��.AA{�	�5�8s�.���a��i�륮`_]Z-`M�%wy�Kck��ݾM�b��R�CW�d�\�\�~ E!���q��]���l5��m��f]ͥ���]����b	�X/vf|֦��`6\���+~/vQnH�M^��gɳ�6�H�	}z�z�=����<�Ost��e	'�@	)�b�g vZ����C�-Ӫ����v��v�i2�@���b����t�o,�7U��׈�)����f��S�c0�6;�s�z�|;��-#83QӋ�-���N�E�w�1���.=F��
���IN�^9�n�%�3�C��nWP�݈��T�x����󌏅�0P�s�N'��݊��3B����Sȣ􂑇@Ϋ��!�mǵ~f�%�\W���?�����#5��2=tR��՗8In�N�B������}�+wq�X���d��`��	�A��=�)��Ȃ� q��IT�Yҩ�4��	Q��e7��w�Wך�1S��XlxVHYEB    edab    1ad0x��&����U�N��0����:S2 @R	j�&���i_:Y�{��Ȏ xL9ݞ����	�P���VK��g�&M��#��k�� 6�a�(O��!��V���Ƅc�Dǯ�����c�K6��H���Y���<��|=��3C���ϊN�#d�S|\���L�'!_{+?TF�)�m8?]�R���0�1���Ï*�"K���	�<m�����p���^�*��\�8�䍧��>�����;'���G�N5��jW�%mŤiG���a�Cˋ��E79p��0��f�)>~�2�͹ʽ�-D�#C&��;~�E~\\Ŷ4���N����!X������r��f��|���!Ԯk����J���;!��Ls�{�����ힴ�7_T�4�P�x P��	
����'O?rJ{<w���k���y��<�7s�c"ٵ�뿼�\�sV`A��6�6!�q�Z�����4]�Q���H3�*�^��)2�
�Tɍt�2
�y�bWi��BC���G0&�k��l�0��Ӈ�2����g������
_��~{��s�'�Gf�:ec�u�2ߘ�.���+�&1�q���b����PG�!��tEai�S�D����3�������Y�6o!L�m�{B1"C��{��In`dTh�R��s=�c���e�ժyCV!/�|�+�4(��.C�q�L ������G�DLM�/�>��pU
�z�l�G( �oD�udI���.�=15Ƅ-��p�����TJ���Z��ѐ��ᢓX.j_��8yMB�VF �5W5��IX˵adg��_�Z,2gNq��~W`���&���Sɐ	ٕ,�������H��
P�~���ޒk߶9B3�1���9��w�j����ߩ�!���T`k^�d��:nE���j����k�#�Mr}����1��� }�=(�jN�5�H�U�	O]?��^��%�.�z���e[�����:c�$ڎ��>&�V�/H�x�"�ݦ�J6!@L{L�r �F�v�f��.nk��b�&��m���΍�^�u�X��3��O��®�J,�.eb��������*���鎳��o{4P�������0����/����ܚ���P��ee�z��R�M\�wQ����.LR6�.r��j�y�\�7�ņ�Tҭu��tB~@=U��t�Z� a{3>��mP�D���H��"�5��U��o��T��8y��Y%��~�ޟ�7o�������R�-c�hT�(���Ѳ%5��G4H�n�5�#�e�<A�!��-u���Ck��A��P_�E���؅�V���e|~�)E���}j�2UP���������c(� #��@��#�~��y�-R�>[�"o:J\�kD�:A��S��;��h������`�������[-f��&e��_c}2���	��ӛ�BO�������W�5MT�D3��)�2�0:8*�+"��bwk/hy�$��/��x'����$P���?e>��YfG� �4�k���b;���5��|���C��֐\3n��4�T	Pz-ɪm�s��o0,,gd���b:��%���T������C�.���6`	�h\"X�2A�'Wېp�>0";�o]"�7<O�4>�v��w������-�}�!,�0�R8#�g쇕�/�?�T�Z����8/�hM  P�M�U��i �c��R�:����@�Qr̫���M9#b7��2�T�I�R�v�'�q�ԋ��2�ż�,��`_������A�13�%O#��}��ETWN���E0�U�������	�w��}w) Ta�;�T����"i��M����4.ߜ���A^�} z{�{�c"jZ���[ Yb �\���|�Ɛ��.5+�4a��%e��8c������b�KEf��ZN�.����C�g���P�6��[9WM���D\ɗ��#��
n�j�F�%3�K͔`�SG��C�EO^�L+�H�8hȈ�';kt�i���M��'�h���O"L�A���[	�����z��,�Pty>IQm�y??�-b�Ƶj��������nw���L
?԰�"�9��=��jh`�Mk�ٽ�G���s�^���;��px�bX��X޼Rf]��ˬ���f��ѥv�%�s�T}jމf	&4�X�UO�^RRgi�lK$�fc�@�E��{��fވ8���u�xcfT���hl@���<����#����R���4�.ϡL���((��J$S�^�%Vt~es@�q�<2>��S����|.Ri��C����S��j+�Ȟ�n[ÿ3b{(�%�Obv"-:��+���RƆߊ�00��G���"-�s?Gj!�&�Q��!������ʪ�2����qJ�dJ�ʿ[����!�a�	*���E�&	�r5lA�>j��o]_C�L�T���X��0=[r��Y�T�Bgg�3���ʔ��'�,!"����D{sZzwa,G�Y
B3oGFҶ��R3\�3D�eo#,�A��~·(��xg�¶�>�C�	8�M��Ħ�����m�$�����n3��ј�w��ЏE������
�vX>?[4)�E�^:�}�3;L��	\lkH�^
��)j��Ll�m7YyW��׈�5ː91!Ԋ�c��m�N��&M+NL�
�o�4,���s�����̸��9g+�W8��s��+�RcZ��=Iү�][� DX>p���%�k�	��e.u|m�=da�����Y�L�#�x��d0���Ƭ~ǥ҉�Ÿ�UɭT� ��|�@�&��ٜ
�>4XT&c���ע�`���S8�Ck9������53�锬l��c��A�|W0޾�I=q��R� �_���.3��÷�!���}}Uh�v��i��?���*y��%�h��Yz�NQ���t�KSu��2�v����r]��l}o�r
T`iR��$Q�8�1���k�`��_�E%@��)�1�<�%��m�Z�Xtmg5ҳ8����V:x�����Q�N�7VEan�W��pl��e�V�Hp��v]���.��'e+�K�^�8l2���/ۭ5����/�+;E�L��сaoU�M-
�a�V��I�#�;�!�7��7k�P1�(P�@ ����c[B���[s·oD����L��Y ��w�b����r 44[!g���j�e]��`�v8Y�jl�$X����F���Er���s�S����+�}������+^�Nߛ�6��L�=��$�ɬ��E2ou� �V.�r�-�R:���&��Q���J���̛;Sư��~k-)L*'>ȏ�x�@~:�帛4�F��wO��C?�1�'��3�<��u����d3�O�'�v�b~��_J�L��ی���Q6WAM�.��w�{���r���Z6!���.��*�C��-w:?c˳����6�M�.Cm~�Ŧ���S c����Y]�#ʛH��(͹�z] \/y(+�Y�U�ؘ�m���t�fL���0�≦yR2�?p�c�f�}�uj]�֤k��V�q���Y9�d��N�UjZH��5��IW�"T�7x��z����:��}���c�p�r�]��GX]�rp�97�ty��00���^6ʻ(ɕg&[��|�_�9�0{�5O>À�t���/�!�vN��}��ؕ�\-x�_p��h݁��'���E�E�s�=�u;Q3WӇѬ����3rJL�Qݣ�	@���^dFR{*��K�8�=�Oz��@�ٿ�	��Zg���I�{T1�w���Z�gt����#;�s?7���9�u�Y&eÜ9��[r�A�'Z����3j�3�
W�������\��P�Lj�=��95)��B~���g�O�Md�>A�f�!Ų���$T�s,:�cbS�'h�8�Y1��1Ð1j�]��(`�됎����(���X��m7��J̸-��JgW_]d*�$?�|��e\��(�k����2�C�=�H=�g���;��.���T����Iz{A������@h�Fs��+b�c��1�m�m %A..\ի>-!`&�W?�(s��y�-�U��}�U:d=�>�\ʺHC�yo	�妋��ͤ ��������� �&������Kn���(Jc2Je}�.)����9k��j�ryD^��f�t��VIY��d���a�k��Щe"[�9��KG?��v��Yٹn�_�H���Tӹ��꣒S�	z����nQ&/Ix��y��*�/��1��8�ux%�-Uq(��e�w�JU�.������Z�l��t��5E3H�=�O<��=#�l(�\N����2!k�[����^}�=|Gy��F�^\�(ʹ1cV*�S�C�$�6e5
�<�u�o�؆�tS껋�$�B������s�W�$��kX��k�j�B�F$��I�,�v���4����3�t�,GJ?�#΁��OӔ����)�(�Ϳ������"���Y����e�����m�c���N:�qZ�,�zj}$IJ�D����?��Z�pm������U\�2�d?�gk��:�/ȏs�P�םl�R$�V�� 5k�m�2����eqNN7���EE�P�@�������N��C�H�*�	�#�ް�	r�D��Զ�cx���8���&�a���av���KX�>�y�LB���H*�~rI�)B� g��,tԒ
�"�!S�4���X˿ь���:�w��/MbS=�����&Dicw���#v|C4�{�+y/��xu�n\�����f{���H�X�}˯M��"�y�v�����H\:�k�ֆRt^z͹]-o��?������u��P�Ee��m�I�K��S�Z���o�GԢ�N}�]�cX����ȩ#b���T�_�r�	Z0 W�z��g��4���Y����b���>��) ��MG��PV���p��v�$�4kN�R,�x6n!7�"EIvm��������aPT�Vz�� �����K�:���٣ҺhEx3	�-8-�!�ji��g�m��)�t���󲗟�����e'�:ڢ�����(>ᡂ�hsh��po�w5/a���T?���Ä+9�x@����T�KH%��%rđ}���|�����伋�:.���&��f*W{Hˬf)���!�8p�����l|\_��A�>.B�Hc�$]�g	�P�
���Ga�ꓯ�@B<[�Ů;͌���
�ڶA��hU����B{�eK��Z�e��ʬsMg�gz^qb{;�G��\�u��M�%-*��0��@<s��vaN«�$�lT<�����tf�F��G��S����x��pV~Z賝�ʞ����/��S���+�.���(`�1��r.Vy@gr�J!�M��d��'�/N�?��#�)���Y`���cE�Y� XPv�?��K���Z,66�	�7:}��MJ&#�(+��a�h��t���;�ʧ�C>�U�E����Y���F ��)#:��#H~�:<
�jQF���F�-N� ��IB��J�$B�ba%_��ǥ!ލ���֫��S��j���9M�1!� fa�6nr��f����a��]|Ds���^h<�8g�d�A��5�]���S�}S��H���_٘�-λ?�/�D�Cu-�s"�Lv�/��vh���{���������
s?��b��ۤ�jM�;����0a����}Zyʟ�-�-�6yu^�����)S]��3�QU]}\��8�7���/��� �#�.i�'�!��6f+�U��}�R��Wx ��x'L��.i�D���r�����|��U����.*E;��"Db5���OS�
�������Co��G�t��N0I�U/�cVO�\�pKH���_��4����V��Y��⻵����_�(�p��=�XJ� ���Y�얎c�03�V���V,����U�ĸz��x���r(�{3l;�h�W~w��Bˋ=!�Q��*��*~\���E"aK���-��w��1,]����k�F
�ҵ�)3��>xx��P`)�:���C�KC���d��O����C��XO�uprٷm��ɭ'��XP�q@�(k����O^H1��*y�2\ Y���J�|ȍ�`e�*܋^���"?�����re��h��4X��$���y�9W�:���g�C�Ȋ17�ﲫ�0�r+)k���l>v_�`���<�_�(��q8��+?�c�N�Əգ��=m<�?\���Еik��G=){���S�S�M��R�J�7���cv�f�o^\#pߊ��w���3�P�$^}k��X|)�ƵOQ���Fl��pvՉ��#CK����%u�S�#�ڑq�b%o`x���v=X@��`�Q;�����]�����V��^A�';��׭�p�g��F��D��v�g�K���t>=A�ͩD;� A]aU�n_Z 1;\�D��Sw���9K�;�MI�_k�*o��Xm=��o
#��k�b�������f~���������(�B��r�N_�Kv�em0X��=��O�ʎ����E�{�e�E����6=�4,h*�B���2@��d�,Lx�G?����-׀��>V4H���:�ɏn0�'�;��T����}^��^��@���j�����Пe�	�Fw���$Y+6��r(�﫻$@8��p�)���⽢���3���2��u[��V���5%���IX��k�?V����'�Fƌl	[�b�,ʄ� J�X������]�7�.����$f�����>d���p�;
`jZQ��+PǷ`��R����3i 8������]%�eb�Y53��n�8���z�IΦ ���