XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��jK.&�h,/Wbh�놂Y��˵��9��0���n�m�pJ�O�I��`��#�]��?�{��#9v�֡��0���H۔
���"�, �Q���Z猞�o�~'4hOf�O!Ţ��ش�h�R�Vy'�OO��-��$����w��>��q�?���-+x�s�w��=[��+��I���@��}c�g7\�l��
-?��K���)w��� %xR�*ÿ|1��܆Pʂl�0BiO��t�� ���%��C/̃D�r0¸��DN��B���@�L����v�����*A�l��#�4]�k��構!��!�8�,_;�`��qsPŖ]R}(f�@}�Mz�pg��l�z.�8-_���Z%˫^f��,G ��kL����ʭ�j\&a8Ч�Gr�ݟP��;��<���B��i��-�"!(�� �>��ꋒ��F�����G!h�}�#2���Ӷ�w��C䆣�٘ �@HoA�V��XIۡ�`����=��"�H|�G.hD�V�-�x�ۋ� @�_k�s� =M�g���	/��z�6���p��Zb�{�V��ħ��@B��ҖU
����ݩ�+�N��͖d�.#�M3��=�*t��S�Sp�Ŝ���RP�I-��i���v�`u�0����65�:��-X`ל�_tEu��\����p��'wU�!n��^w��k��g���Wq.�MR],��	1�h�c��z�{]J�����0^�8)s����(6�UM�=��*�|��a8�؀�=m	�XlxVHYEB    4a98     e80���4GY)3�s�����b�̘��G��b�a����y�U�jf(.�����{'�C�[H�!�Y.g��ޕ1�]H(��ίNI�*��(���W�и���g�<�yCn� I=*f�/4���x��0�(�{�3�,X?�Z6�d�P7�G���V������g4P(k��Hx�x>��Nю��ٮ6R
ѯv�VΫME2�V>d�Ɨ�!9Z7��Zlg���Ԭ3��Y�V|�Gҧ":@��	�z�V$�B��E�C�"������?�m�d���[,�.!1AG6/���X.�9�Z�qrnЙL��;ڼ!�ދ��`7[�q�[>��4����$�'M}"a��uT/����M�;F'�q�R4��E و���N�]�,c��M�_j%&��qul���y@~W)��B$ด�T��]�� ���U�D*(Wn�"��Rx�Ux#���(�s�(`�L2�U�S�p�##zfP%�ƅ�5�&S�j��9޶���e�^	V�n4���2zi�sn�6*��|MF&Q����,��˃n^���a�<L��b��!�9}8��	� W��J!�fmKѩ�=]���Q�5y���Y�� ��x�#�6�ӱ�ނT�nT�����r|��(h`�^@=��=�����vHq��i���g�"aȼ-�'�rq����Ed�]P��N�qY�AМK���T0�� ��Dh�G�F=W�KGot���wQP�9�#�o�x�W ���`V{g�sKo�$?�����Ƥ6�=��P�ƭ�G%~�E��4�!�:O��Vu E�U!��`=FJ����r��C$��H�AFֳF��j2eÝ����V�}���R�G%�O������^2���3��He6�����t-<��ɟhY��(<LH�<�]>J�<;/	��v���/V�i���@V'f����wشtD�7f�������N¿w��Q��4h�@�e�������\��N����x�l��N8e����1{�S�U�i�I��@-����;d��%��ŀ��r��T�����ΰ	<�ԝB��׉/P)����E����4��(,�ߚg@8�W܀ q�Wݪ�M���Le�����P(���
�(G�\����?0Au͆xG��C�0��0tA�t��ŴnB�G�:��ס�>1�R�:��W�60�<�3��X�AJܲ����j	*j����W*�&az-F�R�jFM�bws`�u�6�եx���<$3�l���#9��[���_l]vu<RȄy���ԟ�U]�B(|�]��`^��Ԍ�$ /`Cۙ�:�'T���R`�%�G���'�8�f�w9�A�t}�Upy%�y����Y2�jn@�w(�6�r?��,8��q�a�J����D�'��n�H� {��9a^)��6q\@���/�eP	*�x[�}@��Ԡ?��΅�g(�.!���|X��u$K҈�U�?�л%Ξ�å5o�}��0
�t��Zw� ��R%����5 ����|P�bG�|�G��CGXU	��^F��.�EΜ(�ؐI@sr��U���`Q0F�܎�ߕ�� �F���ʬ7��^IZ�k������<�eG-��K���r�<����0�r�:�m�	�R8��Ӷ�Z���"���NNL�����b�\�𡎷=<n`�"/:r	�.��ٕ����6#���c�o���kأr�g(>XP� f�ڐ��]��g��v-��aes˒{c'I��݉(�ᒝ��	E=5�Atb�:Q��<�Pȟ�S��Ѡ�]�N�����Ң�!��z��H=X����v�'�U�\Pd��
�O�(�䝴���D\F��(=Xb������a
��t�������RE�>��]��S3+�!3d�3�X�Q>����O}J���rbY�+{x�5�����8��W�MJ��E�vg?��6Q4J��elS_ϗA�G�~�JD�$�M��2AG�7�ڇF�?���!��H��&���d�^-@89�'��[�$�TN�o��.$X|���������<:�����q��@���O���])D���@bT�'81�5G��_�.P/���g�: #��~pP�@
�p�T�B��]щ��G�=>#�G��jcZ��L��������掱y{����6H���*���`5��(�àF��S�[;d�9m����t.,��mjB���y?.��
�� ev%,C��X"���ZsS��U����I��iH��g�1+�{�%�v�:0;p;����K��h�<� rv2��e�%#a���w�
C���������B��].'x�Y2�uH����H����~����dp7�ݟ|���?����P�����A�HCb}���Ɨ8e�C�.#��貎�H�0�t���³w�4B�2>C�W�Ϊ%=U6��
���;a�����8T���6/�\� �vY��i�,z@��bU 绿
uE6�X�g��a����Ä��kY@d�2�)U�R��h�e��&T[��;���a���%s������06E�b\>��b|#�B���w�Q�[ftC���dAK]����D��%�U>a��Dq� ;���V.\�c�ה�r�z4S���:[�]���7;(�d�q����p�W�zUn�������r� 6���5��_��Q���Ÿ�ʻ�B�zL+Ih�K�r���/,�����\��x�$u� ���L�Ճp��CPb��~���"��* �4�|�ܶ7�����D�(�_c�Oq��
��
Ld�h�*�$� 1�)��~P��ˍ\o�b"��d���,�ۇN�o��I5�#��N @D+s
$3����uNk/����C���E6o���e���4�4�7IA�:�\<�qL��O��0e��XC�W,]oυ��t9�Đ��RK�H����^����ԋ�����̨��u1""��b���Л�mOل����A`9x�wvuVk�T�2bm4�����Am�,���Z0lۻ��4s?&
S�Q�c�*y96�"V�X!�,��
/�H":�1*���E'<Wfv��[��7Z`X�~Z=#V)����F7�|��`A1�ʒj�=f�pp��f���U��T�!�ҙ�&iD^�-ģP��޷��S��9G����9�6��d$��<�����_����������;�yt����� 6\h�;T���oA\�Q��jl��%�:�W�� ��N"�o�_ˢOH~y܊b4z-i�m2� k����ܬEDb���x��	���s�c� C�ͳ��Ɂ۫��\zB�+_,�SM�]w����Xv�J��N�&�n��k��� ��v��>��4�e�DёG���*c?0�_�Q�Έ�l�`�Ų�v�5�*D�3�5G>Y�ݽ].��s��ٙ�����4��W���g��?U�>e�b�@�*p�}�|h�?ڢY*b*6z,Moll��O�9����9�����p��x^��úv�R��z��<��z"厜��`�OClRv�֙7S8���B䗉:��-�vnS��p��73��
 ���7����)$}���_�E�"-���Ѐ�Z�� �Ob�l�诒x�QU���rh�X��6ܥ�8)+d�;E�L�;�y���C��Wx��=�d�����.42{#��f�Wo����c�i@���F�)V�+��Y�Ap�,`TZ�