XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��+.�kw:��HU
�A�.N��I�Փ\�C!|@��¯L�\J�����������>�DO��k��BM��-Z�׬���>Ǩ���c�s�᱄��4�Q9z��H�/,�-ͽ�l��'����a���Q�j���}{�+ ^�S3�7A�(�����&�?{=jF���CF9T�	*J�<OO�KE�vJBm�,���Ea�J�F��9�#���[z�LR7N��]����c�`xƲ�<�`���uި�M���f��r����/�6�����VDjL2>�CA��{f��#ore��[�NR����=?�Z�A� U��T[��6���҄�{k��[�����*�V��(o�`x�˨�p�,	&�{���Eg�;����9Vc*�|�4dh�h�v��SI� ��IZ�z��2.58Z�(�R�4\�xհ�XlDM�ū�J�!��.�lѷ���)G��/e����ݧN��8EJ�2ԣ{��oy�f���ӎi6��㎡��2�}ʱy��S�%�;�$�ړ�r0�b�������'�T��t�G���L,-&�x���Ip;�6X��2��Ns�H�<���D��'��e�T�0>�e�<�,�%�N�!��-������X?W� ��MZ��?%��`9�x,���:�4"��o0���5�*�D�f���,gtf�nk\m��mv��ۂ��NI��S����f��0u�{7PRY?��U��&aX���:���4-���3w[�>�lȈa3���* �N&��ߠ!�`KC���I�XlxVHYEB    9b67     f50'�ā��Hf%Hha�tZ^�ذ���x^3�2�?ܝ�s�ç�	��ƣ�x��so'�䱒ي�y�KG���ėP�c���`�g�kc��kh%N��i��]&���}���|{�S�#U��	��7���AY��a�!n�w}E��3eԋ�-�U2���8>Y���9j3̷W��C��|�R	>��K�H2���]�I�*k)�.���ᖱH�(��%jG}�=�E},�4�o�z��v�A���QZ�TB�]u���;у�e
���GѶ�^+���k`R	�
Om>���L!R��i�>���Z�
}�ȯG}k�L�|��q� �����*�����Ue<�D�;2�Ǌ���L�ǣ����Qk-&"�e'���*G�ޅԪ<��E��I������_�{�6��&���5��s�{>��$9
Bk<���g�Vǔ�9�0�z(l�`�ޘ�8f�\�Y���;��DDd �q��!v5 ˅���=�eË���P��O�)9���Ǒ<+=8H�r�%T%����g{#��J�A>�T��s*CN젡e��4�L�㗭��p�s��@�Ќ۵k���b���E���a`)����* I��Ӧ�ϙo�����;GT2�tZZ��$���(�Mɨ�����q��ô !+�/o��ύH�
0N��=��8	<{����-3�0��D[�]C�]SKt���πź4]�@˴k�C����˯e��#䕈>O�_��t�4���Ȑg�+�>����"���H
��hٯC�䊑�}V��<�o��H�hG63�KP��U��U��h|p{�YNE���%K����Q�Ďq�wW�d��$[�_�����(�?�u6Crd@�a%C�+Ғ/p)w���$$�">�\�	f�=�����O�]��gQ$��T"��x)T�<���N�Fb��0�iۻ���!�T,oc�YF����6b����bF��/���Y3�h�F�Q���F�c�N� �q��;�-�_��P��x��/~eݚ H�,���}4��$#�y8��F�%����k(3��U�%EJ����jacK{V�������ăU���:� ���:�&Փ�Ȯ�>'9-p0.)��߹�I	�̨�tJ��[Pv���*�;��=���c�'?�]	O���fZ����6�U��I_���z��]N��Ny���̮����!�Yh��N��&
 6=6�Fa%W}4�NLxnY�و��-'��߅+�6UP��ud��7�]n���P�q,��8�A�3��۫H\�~��5�oxw����Qif%�=��TZW�1%�w�9~�d~�S����8uR�ﭥ#��\8n��H`5��xۺ)v�dH}��Әᆙ��_�w̱x	���M����m�0<0ꗨ��W٧�����g	v]��3+)�I�َ+�^@�U&���<�����oJ��rFv4!�UEl;q�A���$�u]��_�f�_����4��:�0yv'�����	�j|�5�S�7�.���&ڪ�
��/��jeM�q��	��K����=�`�cu�gyz����\O�-���ָ<F��>(�+O�׈�U9w�[:�H����!����l�����	��Bv�I��wnZ(O��(��`Bd�=�8����9׀(p�6?z���!i�z_�t'.�C�X����7��q�OP�2��{�X���i����聽��QǖH��;�{5Y�mY;E'(��*@|�R7/,��m��.dn��-����.3��j�?&��*�����z�yq�#w�ʚ��9U�Yw�q��n4`+a1�;�N�'�<�2��76��'���ʴLY:D���.念XGU_�*���9�`o(�fV�< ���[���x��#�A���.�6𘉠h�+��Q&���Y#L�a��������_�p˥Hs3�T��AʃE=A���Ǳ��`WC�ҵ9DS��5{��;������n��k%�:$�-B����C�?��Ԛ��Ԡ�刣d��_�1|��3��G�p�4�u��6�s%���1z�"���ZL�:Mg؝����RD���LD��1H�>�$���f_9��MX���\Y��uR������%�7�*�����9K{��y����>��=��^���;�.SB�V*����l���$7w	eyy|t�=�{^;) �"���S���tl��Y|��PL�g8RW�n6yE� /�#5����z�\�Q3���� IX�3^T@~	��f�(0y-����z�H�z/R�I�� �-.`�A��?Ѵ�����`{�JH�@�a��N�+s����@�n(՗W\f�ڇL���Qt}�Q��I��=&�\����AxȞ�0oi�]��8{�M���`+|���[�b�0)ED_��҈}'��#A�t����	榼R�;�M_A�!�4=��D~C���rO���m�[��@��H�iu�?~����[G�A;�\ nW-ýb?�����Y@DVC����r�N��/�7:�ƫ��g������E�����S�����Fx�H���j֣sO��6�6.�Ù��iY���ʫy?�!o0T��d���e���bJ���MhG]뚧B1%�'w�I��2�8\&
u2C��/�oS/Ǣ#j�M�����T��	;e�g�
��+��<)��@
��.xe����j���Dnx8"p�mW_�t+��E�¡�5��G��D�Ը�w�X��'� ���q�G���MV��ĲF�g]��D�0���>�C��K-LӼi�M��Y=��s�� �^UY/C����~�Y�`*��%Q��]����@XU��5%�v�lH�tg	ʙ��k�å�L�����0�����>fR�<�h�f�f_��Z��[V���q��!�>�B��`N��
�N͕��ڋ�[��e�S�E���t{7SE��!�o��Ɂ�NUs�����7ul�s�)�7cBiHs��wol*HT@��X#��CK0o���-
b��1k�9mb+,�%��(���/�����Ȩ�T�
��8y�1���.������۟�.H$O}���:~��7<�������ű��
�`bx���%N��ܢl�F�@�B~><6�y��90����="�i.��	40"o~R*.����]1��
h���Nq���f��Јc\(�q�_Cхeކ��[O�K��1r��(N��JH�j: �G�,�}�E�O���?��ܵ�$t����ɣ��'6�R=t?R�WM�}��yF��@i�K�&�:#탣$n�A^� �?���s!�/ZGmV7¸^w3X6Bfpu+�o���F��-���
B7���?�8::ʋ[V�+InE10�:�����\}��d 6�s���/ƣ�~MBC��K�Ք���&J6�"0��{�ԣ3���(�?NP��U̘����8�_�rH�Ji*�Ӹ�Sԃ(=���%-F��8���sS�6U�8/ȴ7���1jX��R�U��
#R�ԡ7�]���w���]��Gb�d�/��ݻ�p�h�=� =�g��
�de�(SO(��#ݴ�z2��}-�StR��B��<%h��q�6{`=�{��ϸګ�M�}
o*�����b��]˦J�>��P�͂k�`�Q����;�3���00 >�3�ӉU�8hY���C�>~�|�l��U�9�Og�c�Xf3���D&&���E��u��mjkp���?*e�}x��rGD�O��/o�Z�0�fG�=)\���
� ��[�
Or�kU�;`��Ǡ��`��f����Ŗ�sMB�,+<f��͜S�O�	�<�w�A0�R�����~cQ4��e&�҅��6�dZ¾��	w��7��H+3�_����3���D0�D/�~���PZ�f�{I�F�r.������|p