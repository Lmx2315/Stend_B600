XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���H[/RgP��ۍBý���@�Ԩ/�l&Ʇ�������rejk嘽+�[^�4n̋)*������I�NZݣ)U�V��4\sM�;����ؒW��4a)�kq�+dn,X�,c=��8��v�@��C��.Sn�!bBE�e7P��/6�ظ�S'�g?�*GDzh�_���JKn����8c����<�\ƞ�_�4Q�u1 i��ο6z�޾^)���1zꪑu��sE����h2@�V&�(o�t�DuD�^�a���Zx>���J)_�	,�ɅvE�\�l )C����lfb�+>���n��7��l��16@��o��D��·=���M�V|?�/���ip���.Tl��[e�9�la�> ���?~��v��rdJ���5�́%�QVj��4�6��5�~s�B�J�y�G�M8�u֌��%��zό�;w7�Z`U��?^k�!_Q��=���
���iP ��]ͅ�ǚ~O������@���N�Te�:g�İYcw���*?Z�9N�\�h��f�*��'��HP~ѥ��]j��G2�%�s>PeU��:^]{�`��+�1n��*�bu��'Ū�	����+x�=ұ �6�M��1��ܺ:g��-�B)J�**�M{ƶT��2>_�̘�C�ؔ�4;A	�i����}b�]NL} ���YsW^s�]��S���61�	������w���k�1!)���N.�wm7��snѦ�m�6Gq��eз�榆��K��dY��!�kXlxVHYEB    23f3     910�&J��!]���W�����W����㲯�;�'[@�"͙yJ?�EPK��ݎ?����L� l.�y����L���@��(� R�\G�l��m{f~�6�9zj6��P\ȓ?\�X�ʳ�p�f'ѹ�F)�h���>xi��Mv����Ƹ���x�����at#cك��e�:B���I�Z�q,b��6����2�NT;�џ"J��8���������S�2��P<O&-+	��E���tO!��a���֐��'�X���O�,��!o+�� ���v*����V�-�z[�ɤW�}�&%����ǲӅ��/Ӥ���_\"R�/G;�qw	e���bE��0M�Il���P����Z�/���{\�l�%tF���Å*���'JX�z!����V�{;��%1N�"�;|NAE[��?cE���~I�����揞(���c@NCӡS�DB�(�}��Y�L�%yWg�D�=��B��ȧ��}�x�V�=@����j/\�M6�:�,��z�\B���<��S;G�,@?��`��$�o0�i�&��6�Z=X�߿��7}%�e2��5_G�֯�A͹�?L�	�Z?���:bү���N�k�X�6O��M��ǙŃ$���JC���� �Þc�ګ?�3ãMf��^R�R��7SKQ�D�~�l�HȠI63;k��#�l~�A�u� L͍�P)zP��6=��PW߃���F�G�=�?~l�na�9̜�_!t�@k�]��[��I=�c��=�x��uu,��̽�������������Q`��h/����r��8��p�5�Z�M
.�d�2�Pd��i��^�a��%_�[	�I���{y;n��2|����{踞�;`&&��*�sF�´>u�e&/�3�E\mR������UO�R�b���a�=B���}b��m��(�з�$Rf	�vb�v��k�������g4óbWo]�4 b��1��աꅇ&+_qg��m�c\����ӏO�6E#֡Ag����KI�����t�N!3�,[��(=��\�[N&-n[;0��	��͸	5���� 中>-�6b�>���n��M�^l
 g�)�����O"Q�aF�>��7:�e�,�NI���������\��r��=�f�L�j�}�2�o7�C ��4���}
D庛Kn����i�s��&E��w̓����:�U��UĬH5˩'U�v�A���.��
�\�����q�c~rt\���W���JD_˽�ly�UT�9ȹ��f�j��P߷��
[.�=Æ�#�гT�2DUv}�@����ߝ2v��*��x+�[oB�L�*��&"lK�x���⸁�����z��o⥁b��E����nSja�:�U���oI^�fc���"���0e�f�pG�D怰�5�y�t{�)W��:@r��c��T��S�u��'��s8�׮�x�M�o�1Q�"�S_��f~�I>Se*o �[)�%�g���\2;7�!�@7�Dx)���_8f-�8>*�7��/��_}NmQ�AB�7�7�i�xy��<	?���K�$!�f��J���:�c�pTs��R�~�d�n��Y�+�m�饚pmu��_^h(�P�4"�:˹������uh�U�Ơ�Ĝg�����R*qמ�7��n�	g�$S���l:B=\1��#\k���V���+(�<;����jw$Y�~�������qŋa.Q����~cPt�8��W�M��jm���I�R7�C��]3~�39� ���Д�%H��8���~"�J��],ـ-�h6���
�¦v�8{͖�E���q��#T_X�o�"Lf���D0*���s��������<�	%�?�ˢ�x6���]V ;��q�U�@өK�?j���4���٢L6����z��^r��LE��-�]�������Q ��ﻚ��5AB���I\!Ys�g��on��C��9��NӨ�.{s�����[�#�/�~��(#U���{/!{]$�7s�InX�*WJbT���9,�ɘY��C�7\����@���MP�a�|T��a�Yfr�Q_uT��o�YQ�u��{�N� ��!���w���w֐�X����j��(��e�n`]1�?e(���3��]�q�PMS�fb��Σ3�@xfj���j��v��b��w���,�����],�"q��	�d���V2pŢT1�.�wwb~�˘�>8���ͫ��� f��C�OU�k%8Ս�C}KdʄQ���(Y�]A+��9���v�@��	�E�����"n��/�m߿]�