XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���v#2�i$�)��_�O�_��x�4��^��@��^�m��S�P4��q"����,�d�`Kf�#���)��!j��߱��w�L[����](�p8�6Ճ!P�����O���-�.E�n��r�� �XGU)��r�$&���2��C�e��L���H�	Ϸ�#���;Y1NB��L#a�l�kMɶ-�c'��{В��>�+X�dw�>So��Pn5+�od��!��a�s�^�7��eGNf�����V�l���Jv�7�\�8�YM��=��>+�:��0�.Fa�R�Ϧk�!�ΐU���d�����F<�_���P�"1�K>���Ƙ�(Of�1֗AK�.�X+�$�_w�h���]�pio8i�fU�v>�,�s���ϰyB;H��?� ��]�����</,~�8���Ju�9��n������t�J������Mu\�M��gLx�]���ĸ{М-��m��F��O���v]�B����a��$�a�8�4�*9܅�z%��_
�ӯ?d�X���cFåz�
G��&/��ߕ�f��h��(\���Y�5��0���$c9Q�>,�J�c�����(L��! ݨ�d��j�q�t�<�{̘� RςA� ұ](�C�2��v������Vka��Z�Z�����Y�=S,ˀ��V�o�����E�l�v���j�^�V�j0-���wG&:'P��bM�5�>^�4B��O	�9;A��X����AdS4^O���Q�<�zkY�B/XlxVHYEB     634     250_����S(j�x%a�f|6�]]�����
z'e9�������Y8�/�����,{�6�?�O�k����<�ܕ�mY�V(�"�E-c�Kw~�eE̟���K ���3Y�z����)�UZ�l�$@�s�>qh#��`*���+[�O �zGm]��N��/d����,/9�.i��fL�Dc8V�H��ɹN<�DVE���t ��|������l��[� �έn>�� ���KV��Y�3*b�l�R�U��[�G�8�ӗ�C;�s	��׿[ qXw"u��/��xR	MϠ�}aʆ��^��}K�8�4�����
���ة�4w�������- 6~�e�b&v�����<��13J�8~cv?��	�T*��6fX�M����P��
��W�c~����P#�OK�n�O.�e`Ιȩ�b���Q�QWz��;,	����)�mY�	l�Ϡp��àDI�>(��q\�KC�C��=G(��[�q�>y}T� |�x��_þ��	�sU9>Q��w��nS;���*I*(���L.+-�C�_fX�s�&r<TX���g���xA_��c�*�u�Ѡ��