XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���X���O��f���ȫ���it5OR3��!|L����6����z͙��h?cw\����zU���-|Bt8�I�D�����P�?y��Vc���Q�
,lNL���M
!�C��ه�����+���Js,���أ!j�|r�w�d1+ɖyFR�(��4%6CWG��B`"H�v��Pq�y:�l���:T�>�D��+�����Lw��7��%������V�?������NY1�x�]�(+�zg�pg$+1U)A�߄�!E�9s+��.%���@ջ��Y8c׿�h9P�$�%�l��7������K���1�?#5�$i~�fژv5��qLV��eDD�p�P�20Ua1+���·�Rwo��B�r^Il7�}���U�g�z^�ƀ�ꛜ�1kf�f주ѯdʛ�nT���z�x���i-��ґ�4}�ט��I���i�PZ�5��S@hΏ�� ���]���L?��ھ�;/�%s�l�o7�sc'�L��
�����`�������/�H·�y#R���B;���
���H~\a���b���h��e�� �!5��bVJ��]b&�N����IC�����Dڀ���|>�?^c;x��׿_T����;L���?]��JR���+D�q!\���� ��-���<%�+:�"`x{B�k_��,	!=�t�$Ų|}̾R�ܭm�؞�����Q9��ܦQD���2-��*cx���g��Ԇ���u^P��5�&�/�Pe�h�d|"}<�^AAD"9����zrXlxVHYEB    4b0c     d60�����AEU��=�7(1��A�E�.�Bt$�v����M�R�u,� ��Ջ*�!c-�-Ԕ�U"Ԭ�:Q�'��$��޲�0��B��e��/�Ɇ6}d�cɨ����<�_�$��?�A8��6p�g�"s���b<E�������\��-�TB)�T =���Ό�2�UU���[�����ȹe�D��C��
�� �-W�r"Hv�r�t�4��ں��H&fC��\�턼Ѕ�Qk9�.L�f����q%���X8��q��������R��2e����At܀�_�JVF���Y�*�X_gP�Q^�Is.�c��N�@�8���k��>`����4�,����������tB�KG�M{PD��9,=����^́�ӑn(� �D��W�*���l��z�b*aP[����)ř�v|�,Å
�M�H 4vB�v�CX��jV gm���C�F}#�l,z�Vv��Tܱ�� �)��_[�GT>%!�;�NA�39\�E��eHG^M�<fR����~u6����L/Р��?�飉16�YB�xkU�����e��_��u�1�iԼb���"
^k E�$c�yC�T�����؏QJ[c�=r]��Ǒ-}�Ц�ւ]Pκ�T��y�.8�J���:��	�����L���V����J'��E�sk�;���?�Q�5,�и\�V�������r�U��M�<����`��&��D21�LZ:�APs�7X)��ga3����lI�=�D[�AFu�e_-4�M�}we���S���חt�o�DIVB%�u6SF^v�Q�V�� �sԼ[V��%�u�MC��d�b��\X�^KN}�*e�)6&�s̢��QH�_e��mBA�7cNƐ��ƶ$>W��X�{G�`�6 ���q
�:�R��W+�f�Xd��:^�1[;��,)TR���^x�wA�"StK{T����/)أXT��nI��Byd�|JI��9���U���_�|�*7~Dה�,$�w�21�TQ90j=��ݕf_On6{c/�B
�d��H��ʴWen�Y��Z��4J�Ǆ}ۆ�1��ų�tXDc���|��K����r��)s�|���%�륈�:��������8�OG�`�58ܬ�Ha���b@D~�.�9H	/��D��zDs��&ϼM��V�֛�#�n�8�y[y�Px���咕���P�v���p�� ���GIE�*z��׶��ݰ��O&�Y{��F��U�,�=�xzo�cY'~�a�B���u�@[�	F+��{��8�A�qg���0C��w�oQC@�5�^��ލ�~��^���<~M�W�RŻ����J�5�Q|�&���M,���w��N`3��n��a*ѐ�Nkd���c�UAWTx#������`q;�t����U�L�7S����U�D�������!�Z�&4ZRMߐOK ��}�_<y�hDu	��s����F�9��[�&�`�@Z��������+#�A�c:� nhjf��|v��i��"(��Z�l���>�I.m���Kvݍ��hq����8�{�rFta|���
��t7HV��p�OhN<�6G�����'n��gh^����ьa��r�V|a�ϤnKcjX��f��bυ��б�G�	��=8K�0D����I��Hf�}e���o.��b��C��3�=k@��=���昢���Aa�p��FB����k�"j��+�rcÌ*�F���-�/�%��ŤTB��"�����4�.�:+`JW�f�_bpGm��� օ�7΂�IӚ��)���@3�W�@nf`���ؾ8��#��2�v���y��0i�@��fZUNG���L������}�[JW!�m�����LD~��AQ�!:e��;����zJ>h9Bl	��*2���2�i*�!;��J���΅6�"�ɒ��z烻~��xѲt!2��'x[2�����v�2\���cߚ���1X��h�X+�AP��_��K����]��|�[�H�ji���8r�υ婳)�ۙ?j���&�ֳ�"�C�լ�0��Ϧ� �!�]i=�Q*�Z��	�>#=�V��ƶ���1�]�sU�,�?�R�U�{.�nIā$��~\�'zv,u���?����1B	���՘YE"4?q.��i�~�s����-�\��7�/w�դ���շ�`�2C3���l��R���O�9�����'�-�7+����"RM�3��?
w���'�ͽ���l����ݻ�Ԡ)}tGiRN�SU_.t�v�=�!\~�_P��)����Y�q��zv�#�X��Ø�p�4�Z������8�B��	��<��AԚWҠ���71��{�d6V����D�v���chr��N�j${������(W���7�݅L		F�~�s��X���
rBU!�*|��� �@\& �Y�K`�<
�9%����7jk��/���dv%G@����x]s-�fo{:i���!����<�zw!S:�����`Ҳ?��M���ز��8 �[GUɲ.8$�uѳcs��J�)%M�zU�R����i-O/�Q�g��X��B��:|�Z��rԩ+�e���U!���&Rr7a�^5�	(O��P.���)JF���J8 Y� �<��n�Z �_z��+��L[>D"f�ӦMrM(��k�~15U��-�Q��}��A�p�Tr7w�riE���`d$���N���X"�bD�7�D�whW}��Ѳ3,~1��+���%���M7i6�#��J�S�|�	����tjX��"9�1e�#�
6������v��7�$���Ӈ\�Lvs��\���m�3d���&�{�Y�ɇp��R�,1_�㺁T��.Q�Y���>�rP/�Ƚ��z��*DS�B�%KzQ�-��HZ�@E��R��t��٘�ڎq^8k_���l�9�����E6ًd�Pޭ�3�變>���@C�I%�U�8Y$��V���e�1	"Z?�(p騼�[O��K����#\Z�q�����e3U0	MDl8&g���ꆪP6�Sk��9�8�%;ċ�F��ZCNx�%8��b�$î�+��%O���#76ʽ)5� xP4��X%�K��L{�K�kBo>Ah��5.]*�YL����h��~˞�}x/\����z�������RQ�3�Y�G��I<�祻�<��F.�
�qh���9��?�
�f��/�ƞ�G�4�VG"<X\��*�AC�� 4A�j�(ʣ}�-�U�dʃ�5����D
�fl.���+���jyx?���9yB����ﶸK����p*���X� :�ssN6�&f .NSU3`�K���"�)�I,&���<���iV���Z��,�����D�/_�HQ��SVi8~q�	(�%*b7�_/��>���L o���b3���@������b�bQ��