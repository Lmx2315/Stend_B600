XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��`��U�<#�-��?�4J�ؠ�Ⲍ!U��L�b	{�J`�:ǒc��$��K�_��VuOr-݊e`oV&�-�l�����O���;w-u;s3�l�����|o�`�l7h�칈�����6.�������1�LvO��H�:l�QG�~�M+���"L�gx��ܙ�RP��=���IW*J�Ws�m��|�G~]�3��޼G�1WoE*}��"�����S�i�k"�FV:��/N~�Z�{%� _��;��C�=�kI*�/G�vC�����Τ���a�����Db3��oE$��
@|T-G@�����N����ÇYS\� 3�b�݃��w^)�϶��oc�ԣ��#�~��i� �gI���l:Z+6�
A�z��L��s�6�G:}����p�����l��nm=�r[vJ��\�e�&9DyGRH!��r]U$s��1re�ߙ�Y�&���j� �?p`�vfy⒒�1�P@���চ���k�t6 #�/-9|#���mYCＫ���:�|A#T\�*{�b��ނ#~EMo�]6�����q���=���7Jؐ��3}br�j��,8IOn��[i7��>l��]�|]%:Z�~ƿ���՟�]k�b���>�PO�@�h������}?!<����'c̕}��D��S���@]���<d�!��=h�I߽ʯ�ipW���,��{��9t;�V� w�G�,��&�H��x �&�r���
�M�k���R�+F^v�cY�뜿�Z 2B;/�XlxVHYEB    2861     8d0J^��K�0��SK5�0�@%T�rj�?����������u�A!���T�g(�)N��M����e�E��պL����6�`P���̒�d���j(M����^aq�q���k�;��}tr=�[�Vy�CU��w$�7��L�VZe2�c���{�r���&��+^��� 9��7�k���}Wkx��vo���>|�r_D�B�ɒ��!JU�xU�[tD5H�>%Y�0H,�(LL� ��9�)���y��W�=z$#k�B*+�s�+�� �z�g��i�QU��zA+��
_TӅ5u��vj�R&�S�;`�c����"��t|R/i�z�۸����ސ�d�����7g=�W3��s�LU/��bm|��a���E�I�;�=�>����g��c9<pj�Bq��r�y4X�i(T�ʧ�K驖�����"i~G��)����r=EKEu��B�]����p#;�k�����5�B���hYi��WY|�� ���Pq:83�N刎[CL��ҥ��8��Kex8��>�Xn�����_>;��V?0{�]�;Md�Ax���a[+�Pa��pD�����a
�8]9[�~)�Tl�ks���V7ߪ��-�T�<6Y;w�e6�O�BO$��@496D���6���1Jү|lY�oZ�#7�|Dݲ�!��A.���rF�[*�k&(�*�J3�e��:���h�H
����� $HPx�_7К}�
e���m�(�ؼ�	��(/���p�w��K��G�ncg�x��B�ݭz��f	��������+Wm�/o��1��E�%.`(���'�M}�jqJ��-����.����&D<g����u ,�z���{P��G��x2��Sq+��9�H�KxL;����\K�j���w��ݓ&��ᲕW��_ $��j�	+�:�<SC��c܄D|�:"�̖?�:��!�B!�Aw*�EQ�![˃G�Z�=?�8G��KB3��Ő�?;I�4�H��3K���I�)z68�V!/O��E��@B����_Z�~�$�<�f��3]��,�߯%����$�j�w�#��u�-CI�a!�Q�8K�"��=�i��]�j�;��q�)��Gv�����0�)A�J��RI.��J%>rV����Rы��g�F#Çἢ&�Pf���du$����ķ�i�}�H����5�c����P#�84�l�{_F�Qy`���l��g��Îy�l/�N�VN��sJ������Y�$*&��d��u�鮫��ww��=��~�]RJW�+��
d�H�F�C.�UC�/����U�A��n,`h-�mng�z��!}��o,r�?�܇U̡�n�OXf��H��ޕ̌&+�?�1�_�1��_
nD����6I?����+2~эi�aK3=C�����L�*�f)�t�.C�%D{�֛r,&?LR}�0CLx�Z!G���BI���UU-7ۅ����1(p$�=���h�W*a��w���н�����ȅ��)i�
��eYR����2�ڰ��,TGƛvLʎ�S����O\� [�#���ڬ[����'O��==���h��r�^=4����g*Ĥxۉ��M��+P����Љ�;�.y���r�p���>�nC�x|��0�ɳ��T@��w�a����Ҏ���"���^���>A�4��eZ��qV���c��iނNE����<��$�Dt��	p<���A��V�;R��b𱘖&��0Pr�9�~����s�X�mR1Q���q�7�+#�"����E�at�#�}����,� z��s�]t���<N��}�0�� �֘ʴ�[V	)�,��{[,FS�36��n��N~A&��`�s��K?-6W78�Нēڗm���PEF-��ԄoC�_��6O0c���4~'����6{,�f}�o��L%{~�,����Qc7`2Ǵʵ	��ȓw�{�6�5l҄��듪ML\),����H��k6�������N�8�U�:|o,x6p��6�<M�C�H+���|9���a�RQmCю<�nj��l���Fg/8�3b�a��)z��f)C~~�(SM��S��I��BW�b��e8�c�3��e%m P��an���"���r�,�Ճ�#}�;@+)}&�,�o|Kޑ:
��}1�}6U�\F(B�4�?�GSHǰ�丠$x�lCr��)�x��3'h�XK�jk ��M�3~E�gQ\$�)�