XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���~JP�*΢\���qC�+H��I�TP�n���3�ذF�N掮�� JȺ¢t^��¨譚F�U��f����c����a�S��{���;E?�(�D+������fâ3�v��dP k��oLiY�*��e�mzײ5@��=ٖU:�_" �v�;<iaX�����>�x�(3w� &��E|��'�e}���>���phLbN��ۈ>J��w�����)D����&�3<)I%K �C���� ��dg#��t�\��{��1>4���Z�Rqn��p��U5�p0��6*�^7W���z4��Ԧr&�89yD�w%���ؚ�F��� �d�fh�s��vC�h��i>�&��]_1�?�n�x���h�=���svtH�H�%[�.�l�C��T��� $z[� �H��G��c]m��?�"R�H]�����3/8r׌t��d���C�"�V�I��Q��-zئ
����<�W���q�A��]#)���t�Y�nN��]:G򞈐J��[��z�f�G���﫭b�̑6���&D���7���Q�]b�o�����pr��u�$ݷi�
z��j\�9 $+3�Z���T�6�o�2PbQ�x|:�HG��K�����:��C��K���/M)M��[>����ǃ�d�W�H�~y�Ъ �$2UЩp��vD�\�S����J":l���IhP�Q3کU�]�%1���3� �+����ǹ�\��v��Bx�"ۀ��H ��7C�Ow�+���U$�XlxVHYEB    b892    1b20��,'�b��`�Q���G��d,{�F��;c�Su�p��T�M��Ê�2ˎ�(�twD4Sf04�!�A���TJ�0АL
NO��f��ﲗ���pL�)�R����������]y0���v��P�~T������?q��~��nH�CMj�g^F�$��r� �bO���U� �Ytf繟�Jj'p��i���2�)Xf�#����ڼ��@_!���l�#z�+_D�S�ox��D?�	�h�(Y#US�ӫ�2zq�d��q�g�p��m �n�j�A���[H�4;O�w��M�~j����(ʈ@��1��hY�q��j���-�X�6����]�w���L(��������(��͕|[ �Å C���c7f���<I� ��D@��h���ju��o�B]տ���G1-�q��S�w������t�Җ�+�l)���ͣ�\��6��P���RsBE�@d����� ���&U����;�
1��V���B54A��nR�\vf�!#n?��0>��6!�l����.���*���A* +0b�=*k hˋۂ��;�%���	dg��|��R�[���hg�%�90�B�Ň�tP���j��?�H�/�0��]A�D�אQ��U������WqvBuF��*�����j�e�ǁ�%dN���ÙEr�_��b7"vO�gl>���Sw�+�	��O�V.i(�׼Ϲ���;2 �Ƚ�U�O�p4�d;N���|��y��{�2���oo�?�����\�`��[�]�$X��8궴CL�綜�@W�X�y�7��֩p��f#F�k._�Lg,�o�!n����rÇ�:.d�̕������a�M���Y)ڈ�ٞ�ta�N���؅/?+/S���.��H���	*a�o&��ga���t�X@��=F�s�q��o@Y$�n����PP*�#��j0�PX\T�+���{�ܵ�޹�������T�|1��-�a���bz�
7�j1��0��0j7�o)�� �
S�c��s���'3j�D,R֪���_?�]����I�#r��s��Ɓ�ze>����Zo��[,���6�d�!@���xk+��d������h�uvM\I�C+k�\�E2,lSi��|�ko�|�h`�S�&� C�s$$���1=�W+�͑\ �<k���@�ofl@§7Z��De���_�����:��g����,N��H]�h�����e.�c1wsF= Zi�ʮ��s���rI,����r���p�E,[�,L�=-��������{�����a`�d̈́d@���w�W��+
nRҍ\������
G��5�L��D	,o8�F�o9�?tԻ\^�`��Hm��2\!
�]R'D�90c�e��i3�
�2_���.��TչFX�v����i`������\����Kܩb�jG�����at�Q�lR��-G���Zt0�O���6��޾M2�%�*�l[:F �F�Sv��Pz�x;I��W5�#�|����dZԟdHN������`�k��zmkP����=oA{���>r	�YW:��.�`�d� m�8��A�4r�j�$�rD�լ�JI������;�a��c�
y��i':����*i������{�>���Ă�Qo�t�j~�x�v����!gvlg@���5�g��pg�y�+�Θm����	��_"���r�/K9%�r1���3dn^���-�RF����I l��&\-�������1#u�s�">��:Տd�O�rX2�ײ ��p��t��v//�K+>�%(EѰ�ͽtQ����\	\��y���#	����@*���p�]��ذ>4,�
mϤ{K��u�X����2��I��*����4N)R�7A��D�2��eP��9p��ڔn~����"�A	���ʜ%��|�����8"`#U�a�F��1��<W,��aBIYħ�}�������O��}¸�������W֓c����?��;5>�Pc�7}����|���=7U���]�����,5�eQ�B"Ü,,��v��j���Ǐ�%X�����6H�PE�!)=�o�Ѻ��W�!ȱ�J�~�V�*��n��� ����(��}��[K�U�kV �z&}�0����m�b��R0�r��@�md��^�����;����j�<�n���*j<z����>%�9P������#ShH��-\1��\5�pE9�%��vw�A�!>_�6	)T+ۚ��_m��I��El��\}��t�?_�����kX)���yI�)$f�b5If5�7x5R.�����e�CP�������=�	{� kN܁]&�e�
�@�q���__��%������\S��#��o��p3�a���H2�f��tnFQ;��Rk��CB��ݷ�jC���=Iu�.u�*���X]Y��8�.�w���e/��(#�I��}�%$�p���ة�ȷ��H_����.M0�6{��l��c�[��y��rb���2�l�$��b��/���"q~J0I�cM�&X�+f�R��'"ݢ`��q�MT�$a@����{����H��r9��@�K���(�[��s�xX�>pNc�]�Q�b��8/��=C�z����Ne�	�h�+aD������\G)�����w����l�_���3ex|�'m`�t��O=��bK�����а�y�0b�l�>���*�h$���F��wf�|+�h6��1�e-{��A;�������ڀ8�Zy�����Ef�;�Ի�V"WJ9�C��9@��
�?ig���p�R�%�U,AO��]L��ݿ�xD�����!nG�>�<�;���t��@E���Ɇ�~	˳e3�	���ᾢ���S*�-���A;�=����^���E�x2~�"�tӊu��}�Z_fd����k4��>|.����v�yU���O��>!ߺz{+��)���0˗�0���3�ɂ{�?�[\5!]`=3�����(,Ҽ��j6Զ��^�e�F&�xÄ�5���{JD0��z��%��Zez½ߥܑ��沱P%�ϓTc�Q>�U8��d��(�:�"�>K��e�+��%tLh��ؿ��f��!?�Q����Y����b:E���><�>�[�3Q�c�����*��k*���df5>-�nc�0�LX�|Ց�i�	M�a��\*�Y��
������_�T�V�;6a�5˿�%Y����LA�b���AXS��Yj.9M�;�,�3���ʭK|HTӱ|��9���Ĳ��J8��c� i�K>y]��S��Ó�B�6���?����	t� I>�r�,�Ʒ�K6�B���i9S�q?��P��0:���6��ą^Ƥ�׍ct��$�1{e+7^_����pN�rCB`"M��  |��C�p4	L�`����ۨ���s�%��,�O��"� E2Mr��P�I���(��u��{o?6��w����H�? �����0X�%)�V��=�p���(���-6���6DمX����8���#ъ�EHFl۝T���H!S�"��M�I�8�װ̧���}����ڠvt>�)i��$�|��w#�-|�1�����8#Z��
�>gP�b���l�O_�m*��1�4���AsT,��h�l�t�̫��ڢ+$gwZ�a-����"#���YyQ����ǉ��(([� �x��6�1M}s����/7�|@�2|Lm�)x=w�+s�$a�}F�{�I\��.A���g:�U,զ�jaa�y����EU{��q�6�&�8{�j��V��H�UEY�(*���iC!r�hI;��T9=ϫ��
���17�G�ۨ������F<��`����Ϙ����p��o�����<����񑎖�3��7WMW侥��A�kc��LV'�ޞ:�T=G
� ^q��#�>�Ct^����u\��<���.�?���em�l�#{y��8�Q�r��qM�SA�9�K�����	G�w0u�Cb�G�?�n(�@������n���r�?z1"�vF]�;�ؕ<tU�Vd,Wާ*.ء"�6�b�_w�a�Z�I� H{�@��޺��~ћ��[�d=�uUÈ9��Q
=�Q�����{ ����#N�)�?$��2���E�ӗ��oʱ��i,1�!�,q�$D+�t��ɻuS��زh�ٺ��k���׾�G2T� τu>��l/�6ds�m����K7��9���un�;)؜���R���9��6E0�M�����[���D�'|40b7�}�GS9���5K]Hm��������Ĳ�<H
u��N@�l��D�8��}�� s��Hyp��ҥ�ͩ�I�.~�]R��t�ea`�M}�ci;�C���d����6{�`��y�:�N8KF�(?Z
m/�\0D�w�h��Na��Vv��'�[�7�y���K�Y����T�_f_�� }˖�>�h�F�9�!�e+4:�I�x�h=�,YF�1�ؗl�+j2N�-�l}�i�Qq�(v����=,���8�9�|o��=ȕ<�2\Pq����$C ����T�]�0
"�ﯬ���g��p��1�����Jm"�%)\[~�YV��ib~&(�>V���cb�y�K��|�8����5��ݯpƬi�<)�c�Mͬ��xK��M}j߭�\����We�7M.�D���R��	3�L�?��
�4�1f6>�.��G\��(b�J��w�42����C5�B��.�W@&w�t��x*��U9�'*�0��8�K���x��	�1�����42ݍ[f�dOQ&M�MZ�F�����1<�!A2!���m���Z�$�+�vħ=�4�u9�1���{�#s:�<���3x�N��I؊Ԋ.�G}T���ͺ6I�i��s��T��D%Lќ!��b�h|L���<�#	ȹ�S�H�$�\9S`����KJy��+SRË�v��}k�?���T5�>>U�	dR�M��TN��iw��b�1��	$V9��<�e��{�SKY�g�G���\,8���#���M��f��8É_H��#���PQ�*��؏?�Y�J�&�͂L9W+6CH��vEF"���^N�7Ge���#S�%�K�I�)�V���W���:`�P;˻h����q��%�����ҫ1�Fn�<���/VTǣ�8�\@����>�|�j�d�E9�M�TW�ռz<֧٠��a��F�&�;]��l����Rs�Fcu���+�#Bm����D����F;$1k��e��V�I��,B>���F(�O��\`��r7�X|��D�fWҩ;2���RM%>/���.:9e����q�#���v�Q�-.��x|���N,D;�#��қ����ʔ�iՎTk����drI5���#�Ї˘^ӽL�|�Et�7�M��C4�8��>)�&�W�H�9����;�E��� ���O�@kş�IQ94�'���b�;q2ekX�И�ڦ&<	:V�I[�Z��2�1\zb�٥����t����/���G�`/ ������ŧi������tr鞕Mţ�����M�n�n�/�d�iX�,,L����V)T5/��s���ՐC:5�Տ�D��iDJ���$��v�.�N1�=R 6�'ʽ8�"���#؁_}Z�:��i
.&kx|��վ�xϏ�][��$���KU7�󣖝�)ɽh��R�q��f�e������������T<�^M �yO���{|���꩕���t��.�R�@��l���.����#�Ӓ�6`L�e'i.>;㣙�_�P���L0�F�5�H&S*y}=���>����s��.��	�h���6w�)��_��n���K܀ߚ� ��`Z����K�]yuX�ef���Ll˱4pBs���ۛG-�n�@���7_͟
=-V t��O�ϲ��`^�Q�����2��l�~�����3�XK��x����!2����������7�O,��p�Ă^�J����`��[:%�Ǵ/:�z��ȡ�}���^ E�\%ȇ�����/�ي�����,9�[����y"��(�BR��D)��UmY��ɽ|��?~i@�#�1"�:��l'�>�z���^W�^J��ξ��Z��������>ypY�.� �N���2���~̫Ra{��c��#V���l��klA{��
�`Ck�)<�Y��8;d�yE,9ք^�6���������?��ZqQ�nLv*~��SP�Q�d<��G�$��_��A"��������џ�<�\tF�Z\ޣ���֠n��ci�����5T���w�Y��824QT��+dSv}`ڻ���MS%�0%����Ջ S���t�]�^# ��q��(�L������Y.,��3Ĉ<A^Ǡg1�rIY�C~�jL~&	�<����
�/&�V��c��zQ?��Ձ��<"�o��Y��=�6�);}�54:#����Aw����rG����O�*hwy�}ʄ��=��A�0"��z�ol��c�o��v}9]�|�5-��:��(��`n�ȼ�Z�oi�cſ�vr�+��Š҄m�dw9f��}�;��ur�?�Dh��V����Fx� �Q� s ^����'(ec�>P�Kqٞ3�!�Z��|����CfT����B��C.>�\��eQ���Q�+���Z��!aUx�$
]}��ϻ<��o�ʯ�n��ŏ�pż����d����G�v3o@.��ۺ�,R�
o3B2�#f����a���bz�+��u��z���Ŕ�:WY��M8:0��+}R�ƢM���F,q)�l��Q���ȖG�"?���Q)--4zo_��.�G� �Q#SQ|�	��
oӨ�OxkO��������1�EB�M/���`�h�l��e�L/u�t<LA����=n��