XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��^7@�9GErP��d|�z���U�Y^�h6V��@ݘ��X�*�����C2z�0œy7n(#���0J��LZ(;.��/	�0��;,��["Z.�gO�P�iw8 �%r�|�Ά�H�*Rh�姉O/DۏXĪ�+�a����ג6����q;T;���a��1^;�����^8�@��*�m����؂��cPw�-:N`���䕖�"3
8O���p^!� �B��},�⏁U��dYR���;0�~�g�r���n���T�|DF�K�&������<@��%D�Wg��KR~���_���j�J��p�j*�^d0���k�����s�h�O}@!�i�3i�a�lK�l~���	�ؿ��t��c�(��ڃ7�𾃳�@���]����l�[+�~�e�t��]�u��K� ��Z��X��H�oo�'8ޏZ?Z�%h�jp?4r���H��?/~�;=Č��2h���U��G%��I�2���	�B�B��ZL�;��@�6��چG�I�O����⋪l�1<��'�!%�Ap<��,d�g���B��Mw�?�i��� ���B
.[�'%<��3�v���{цv��OH�=orO��L�p�7��"��K���[ ��~8R����w�-v�}�V�� ���\�b�E��/(s��n��sZ�e��n�޻����]��f�,����w�4[�����bAqD��]d,^��(g�����@V���Y�����E���IAfNp�y3^y|[ܮ.XlxVHYEB    6faf     c30by��s����5wց��B����$��ąO:Ap���԰`�DjY�"2�[�'�fD��x:�����u����nF�٘`|����Յ��� z��CA��s9 ne<h������8��v�]�L�
�菑8v�s�[���>�+{0�&�BI���-{����/� �$��h���t���D��k����yo�Z��2�a	�W�[_T�2˰�>8�遆tlX����:џ�a.y��Mt�@�$G>u	��X��/�Y�GS3uVWc�o�Q<����T��m��G�Ĝ����tf���s�7��G�u�'l��� ��*���AZˆ�A���&�`J��Y ���"�C ���o��W��^`UK�*��Y3�W��0h����6z6�����솱����U�V����)<��Xz����z���
}�r�ٙJ�s8`O�-{#�����θ������wȹ�$�`i��D���C���AN��dj�>��W3��F�i������&�'��0V��+������$j\֡��m@���Hö�(q�	9"s��ʟ@���JUǄ�m�X�>����-���S�Ty���?8�%C�U)>�G��Ӣ�a�Q�ܐ!jW����j�V�ɐo4K���vb,2�:W� ;nsvgS����#V�rGxs����C'J�P��q`��i&)"��8 ^��:/��ť
e(J�Ͻ+�}PB��&I%��4h�dUU,u���m#p��O
����_��D�/�.R ֶ]�N�4�� ��1Xﳫ|���&��M��cy����.a�_���!��|�XΣ&'6�1���.r��q���� Ota�A;��9��+6�ӱ_�X����V�*��	)E� ;�E��;������R��	~{�`^�(��?(�I>�b��@�+��S
����-dAvu���S*F@�bbK�m�6/=��,�v8\R�D�g����y�w��2S�naJ��t͵�����OSE]ĝ��f�~R;�o.n��6=�lgp���7ʟ�Uf>�q̓uV�m��(xqKw�u�D�@�/O1:r�b������,YHږ���8Q_�&�̖���؇b��7�߈��0IEׄ�}!8�#|�%�k�I�7�_,�@��\����b��:�iF�Q�[p�:�l����@��0ڙ�w�в\���x���s�@lO����K�2H�㻷I�_�n��&=�C���O�����5�T���)��_]��~3�����(ZG�MK/���y0�<�i���[Mr\�3�N�`x�fiW4��Jn�F6�?��|{ŗmr�F>q�I��
d��g���ܻ6 K�KP��������u.�U�ߪ��9K�?SX�=ln��J��@k\8.�d�Dv�~|���e�	���m_|���U���(���b�ݔ�/���g��v*���S3t&:䦵M+>;���<s�Ho��_�ݰ�k�f�׼���T[<y���=w-v��5A���_f�!��y�2����n��s���*�e^D?=�)�`i'|��a�L<7d���u5w=��Q~7�]T�v��'��Qʪ���T�$���� @��%W��6Iʆh��=j-l?�|���Dx`�%R`��h��.V��+� 6O�������Dn�����d�L�\��j���Y��g�'Uh��N, ����/,B	�*���A�	_B���H��<�8L:.��Z�;_%cI�j5cA+���<����c��8�-� ��T���[�&�.
�ZC��ʕᡏ�a��T���	�4cߊ_^�����R0u�u�?���!��l����*b��!!�������,�8����V��l����Rl.u�Ews3+:�V�5��V��M����T�|Z�*�N�Ӄ@M�w�}q��4�P�� ��	~�;ʽܜn��0��h"z�t�L���Bs���Pd"\��'���(I������pf��`g�*}~�2�]��y!3�ss���ܾK8ͅ����*T�#E����Y���A-5��d�P�*���e�o��|�GS�c����*�FG��Ͳ�Pv<��>���o����IqR���w�������i������k���f�RYK��:m>(e�`O&�ҿ�F�E���Y}S,�2Կu_1��.�&��ɐJNo�I��f!4Voe"I���NO��@�[�l��5^ا]��P`�c�Rg�z�P�Qd���e��^��������hE3���"�T�Bc��+��!�	u�}�IԜ�r��2p5.��3���]�N�\��U k���K¾y��r`[*9�4FȤ��$��Cd	�܉���[(U8���yC�>064�1��8�
w"{���v�|%x�'�KUQ��:�1�g��]D��_[��΂,��t:�zx8�O$�Ck`f���
P����p1n��nbh��C��̒Ƞ���v�N���H9��eh���S ��R�w�R��l�T� �Kk���]�)�|��q{�,#������+f/�λߴַ@�k_�`�z�� �����9�	���i�Ӡ6�W	���=��\v�?����Ǩs�y�r\�b`Thw��a����)'l-��zfЙ�Sf�Q'x�f�mSF�9��t34��bcvT�vUTw�m��xha<I5���䘟0E-���m�|���}y�J5ÍC���O�⋄�(�����à:�+�75�;3��$>E����oZ�SMZ��P�gYD�'�+�j��F�?�|Wst3����!xȗ���GQ�Vd��-��V�d��v>��H���|�C@,��#w32�q����T����e)�!�0����F����xp"���C�5�^ԓ�$YBKKq����+��:k�]_zSnT�*Xѡ�%��R�Q���T�s�(�B?ᢁ~�,����(�j ٣�'S��o{��(ꪵo�02"��Aޥ��k�9���	��^E	�1a�今��r4���V���SnЮvO�&K����r;[�{�<��j^�Q,`9��8�:9^n���PǛ������/��~=�M_��B@h���̩��5I�h�����(WS|��UM�+}