XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���{���\a�����D�zK�&���O;U:��hN86}���8;8��;�u.��^���to�,UC���f��q.@�I�`4�� ѴC�80J�c�Ɣ?� }fU�㎂'�G�P�;c�B~Y���~�IbbU�2�z5���r�O�_��g��+w���Y����Tꏓ?�Ob7��p���]#�<�v�1�b�-��LAg����7~h9��ߙd7�zw��'î�'XZex?�P��	tM�6B$�!�:�HGt�q)�
.���CE�ૢ3󋃀�_T��/�<���DJ �E=����"xtT��7���4En29�cc8Cg_��'��t:���m���ܑrĠ������\�EZ�[-��diDV>[���^w����ͽ�!6Q��wQWo��P�������|e꽬w���F�*��L���u�� td��������Sᙀ\ѫ(������Æ#���FCz(n�i���:`�X�`ﳏ
��2`�?y�D���%�(�e��NxD�aγ�!�qMJ�;␘�.� �s��Ǿ���/��g�2����6�oä�[i/
r�Q8��η��&��iy����Ы.��=�D����%���GE�)>G�p����G���]��p���~�(��x��;D��	�������+�֬�kP���"~i��^�K�"�H�Ult��:�}����z8�����W�p�(X�^�J`��$G�r3-f�l����r�H�<����Hnb��*�R3Ʈ��G\�.N�XlxVHYEB    a354    1890ԑ���1�<,�|�U��t#p�R��U����+vvU['�9����������Zp*;�P��_K�"A�C�	�c9l�����U�)-;@)��؇��/�ДK�>8��8����
?z�[k��Q���2}�jЖ��`��&g��p��^��|���+5���i:�ƻ�Y�%��'� r�H����_�p��3�Ѽ���0z 9~m4��>���X:a ~p-����;�6 �w�F��>{�^r�9��:K�����B�[���	�Tj)h��װ�8f�Ƅf��O�r���ߝ�CN�l����
9�
8�'��lTxd�ҲN�x��xΌ,}�^0������^�툠J��=P���S���,,3L����88��] c �X�y�4m$���3��4h�������a���(
���Fƍ5qR| �b�����y��r�h kٸ�Os_"�L�K~���]�JnW���M�m��o�tB��£�*o�C���N�pe�7��)(��- �諠(t�֤��{����b�dJ+e�h��Ⱦ9��tx`�^�ٹ�A�p�hyp����S���k	�
��T��ԹqFw�$܁h���]�bϰ� ���Z����0��9���U#�||�/�y�,����7�()��]_��ZR��=֤ː�<ar��h
�}^�w�=+:W�WT�b?s�K�o��{�L��vd���V]�pI�EI*��I����P�Tt�C���U*��*&��zW��.�i�@R����MXB�-�S!?����2��*���u��j�~��N%��'A�y��$����@d���t^�9��������I�YS1�=����o��W�ÎR���&x
�����N�X��ޝB����^k�9��X_���s�.�3��@p�<���dWj1��^n1��Sh��FM,}n��B���4.�\d���ڽ�BBO�L��/Ŝ�ɣ]zU�M��8�@+�ֱ~���"�m(f� F�1Rz��(��?�wY�h�u4����>��~4�	6'��kHT�v�;t-�<����+��q�H�N���soDO�J��H�p�s�5����>$-Z��]���N��B��z���w"��^\(	�MY��b�X���r��.Q��#)�2����d� s{��(-jy��/-��H܉ϰ�z�.wܵj� ��	���.$#�N����a���sJ��Ku���G�ڥ����v�D��HM�z:v3�T$6��#��S˩��z���p��B/p���L�2ӅTڤ�?��9����x��i��H�=E?�U�|���~8o�Bޗ�K-&>{B�"P���1����
x�n-��{�I-I�����tPp)�5 {*��fM�|@�u�����r�m�ȉ����Б�����D]��N` �\���U�y��I�V7���Dby�*�G@h���ivr�s��"�7d}�m��nf�����=T�Xy;X��5\~�+<I��^�}K�"J�1��ŭt7iv�ÉN�\�� n1>hGo0��b�x���L]+r���@�X�`��ʔ���E� @�v�]�ag���,��&!������Y�!غ��.�`�:%��B�1���a�(V_����K��=�Lm��!H����j�	�_>�Du�he_<�`@.q��.�����U4l{� ��%7�)����([��؎v��Ml�C>�FaW��'R���X��-H�����v{J=/WQ�NZ���ƾ�<��0����ͺz�)<�3}/�m�ERap�?�aZ&@���go�><`���=�3���rP����1	��z%�*G��s�j���|�]��9�B)y��RYx�/��~9���:,��ܤ��-~�0�nwxM(W��3�m���	-i-q�0k�1iJ�>��I���DZ�� IF�}�@�BtHWhXld �tT:E ��37�$M����`�jH ��^é��b����2F����P�_YGd��,��aW���&�L�A�`��<�1Nr���	5d��	|�0m׍XH�c#����|Z��X���B@��_7+o��x,i�`����AЯt҇��4za��W��w<ܟR�#�c��J�m�I�(FY,G[l��oA�<��cUov�^e��+�(�>Q�D]Ԝ��&""�*�������y���`����d�|����Vd�("�A�[�BB���N� �J�P�1��&�w���mL}�
轀љ��M�$G��t����e�J_�'���z�Z���!}aJ���	�l#U���p[v!1�����ăK�u8���T;�l��|���gV�/]��)=o0�1�Qt�f�1��e�͕��(N��ϯœ72�Έu��ی^�s��x�.�vw��2YjƓ�(Q�,���&Zk1���e�e,�KV�O������H{vh�s� Q��ctHf6,.P1!V�=r�P�!bcO�������p?z��*�+:�7��i� @xc��Ǩ�kG�
t�QR0H/�5D����կ�D��r�+�t���y������z�l����]ԧ ��ݕ+"Sr���{R��X��r���h�iI&���r?��M9[Hv��i��5�IW1w^���χ���7�N�Np�p�6��J�]#�}��RH�x~aW�)\6�t��d=!����q&¸Rhu����!�X��"�5R	a��(
���[Tt�ǫu�M>�g9�g��D�l��0�萑ќ��	��;Y���E�Q���z�hCt"s���K��Ix��矺eY���0hԨ��2��	FG��%����|`�lի�[F0��1��b�j�'���7���Em"&��!�V���������s�<
�cT�i"c&�w<�b`F��1L�,��V�B���a'Do��81�Cr戈(@���{����{A�7�[�]"��ɥ3�⧵έ����p�����di��@�_��y:���eGZ�B;B���<i���2V��M��z%"���C����e��y��/���׋o����*6M�	��0�[-(Ȱ"#��X�e��u��xs齅E
���?M;+�驔�������[	W�w�8��&3�	�t2;��y��.�*x�������:�����ԩK�ׯ�B�n�>��T���=?��Y�ei9�֡�$c�6�gvj�G�#����ǳ}S*	D�x{}��/~����n k�,�tS�L�I��c�@�f;�I�'AҀ�� q��.�T-A�[*��5f�w7vc�4A`#(�8����M�
u1���`I#�����V����ag�z��G���d�}�"ruj`�H�9�bѻIK���<{z�32�{���q�^;H�|fɷ����\�9�G��E���DY���H��]3������4���;1A�������lyF��� c�J���,)���%R�%�{���R�*�����C4~�:��j U��Mݎ��u_�=q�Ar����͝�آ��7YM�5�{m�x�Q��.���k!0<��|�O�(2��1�@��ɦzj}&0��J���9>wq����s|X6~%V����sb�p�����Lw\M
��i��������m�~�g&E����#�i��+��c���b\ lo�R����J*�@�T8��*s���S�X��BOU������l�X�O6��6���_�G�1�%�H��K����ϟu��J6�xl��>-�-� ͛n=g�Wd�b�&�a�c�'_@U�K���n��P�~�p'F��}|7���O�6etO�M'�ȁ04�H��9���#Ǯ��A�O2�o.�t���Zi�"��\��M�z���m-0c�8�&j�eǸ9iI�q�o,���VQ��y��2��R�֌���zr�ԭe g@i���k��)k�9 eII�@��D U�J_
l���RAwȵ,�	Z�L�<b�4(�u�P��e&zH_A G��"폇��������nϰ<��fM��y��<Y"ot��Blotÿ��Qѵ�֗>�21�G*��gE�_��fF�v��	BL��Z;�+z氻Աkv-)ހ��������_I�@�)%�Z�nz�!�s�{t�8�-~���&ͦр��O��ֈ0_rS�Q�$���7Ϲ=u �;4b�#Ho����Qq�Dh,g�1����h�0?*�X�A�4���X\�W���yǥ�����58͟�V�L~IN���`����$e�ͭ���e�'�;ZPzv�n=�^)� P�%9�d
� ��E�f��5��<o�H8��Qp~mJ(^m�)`
4���@p�j��{���N��1Mn�{������R$Vqh��""[���~�h঳�ZOq���}g���|$���������:��V�O>�`	C�T=��"� ����ض�v^>��'���[٭d�����%�d-4�Jl�O�fy�?쬜e��?
6�Z�n�̤H�G�d3�i�����A
#���,�@���D>̕��v��u�{h�z�eF�VԐ�	�w�:בFP�E%��M�#�i���;�P�\��||Raw��h�f�P�gͪ�	B�e���d&�ow��*�=~ĒgPV�����HLa���ZtΝV	�T)�����MO	�;�9�ph.�ŭW�P�]V�뜂��5u�N�K��ͷz�$��B����,^�q^0�	��g������U��	#/P�77c��~�ŋ����q�8��+Ҿa<jl�Q�o�d�ϕ&;S͜A��F�V0U]v�)�{��x~K-Q��^����$U���ΪXRFbݦ�{�~�H���@�=�-�v
��'�z�o�$�һ��x,Ȧ�i�t��Ta�3E/��3az��%�D��*�ϴ��n���×�?ްZ�\e���踭�n3� 
�}�"�R�o��z�h�i-YNy�C���8���pN���4s\q�/k:�rRL-ؘ	u�M�gL���L@V	E�WP��N)O�����?��暴�=)�B6.'��^@Y�fQV��6��h^�l������0D~�������\������0�o]��9Ku���sz$p�zj����տ�{�7�ٴp�=��B�������K������v���O	N�r8s����/҃f|ؕ�����Τ�n�	a-���h`��=���+S� N����fE����	6��\dYJ��rl�twc�F����n'���#�鏮
��������s��n� ��I�Q������UK �9̑�������=��;
����F�Sz�ɡ���[���dg
��`�������Ӥn�};���� �^*C)��܎a~fqN[��.��P������,E�&�9�Q����Ӆ��%�``���N�A?���y���ئ_h�)q��������3�w�+ܢ�G����v޹Z�}�����8�Fs�&�y�P�&��/V���<ɡ�ݾ�¢��c��"K���z�`��{�i[u�zՐ�6}G�ъj3o<�M��\�-HRBw�uP���D�ɔ���/�P���þ�Yk���L�f�94g�a�����D+'�C��~��0e:͹2���c╹ɞ~�ec�iD�{
ҾB@�7/��)�Ϻk7Fo�Bi�=꓊�I�M�#��s���e��Z�@�"1f���tbnjr�Ǹf��vเ��3��t�@�O+S𝯮�)9!��T��	q&�ȩ�%�����������=0���������Y�>�F�fK���*D!L��:�Ct'�LO�<�r-����!�����,�h��櫢�a7��#e+�E���FV�ȥC~Wc��x���A �u�]My���9����u�8��/��i]&�:X4����1���{����W��)��婒�S?��M H��K�D]��Ər��v�� P�-2T�� ���ouѨxGØ"���3��b?3��*�:���)�^;�O�c�KS�8����歷kR		��׵����// �"�D�@���OH
|���vf�":��Sz�zl�_���#���c	�*ڏi�Ln�s�\��V1ۖLX�)���R�ROq{rȖJ�߅���D�W�VaT�N B@lr�bįސ#@ǲ�`j&j�}M�	��+L����	Z�	K�@����0҂�u��4��	�JV-����90ҶMԢJ�f���̡˿ˊ7fY�bgZ\��R�,�j:�`��p2�2�$j{iV{IOS�|�y�O�eJ�Iř v}���=o�cT�O��