XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��՜���픵:��$�,y��J�p�T	�ݓ(K����b=+�fk��W÷kȤZ����7��V�G^I�����Ԏ?��B�s{���@a	�vs����z2�����_�f�G|Y�頋G^7��]�w�Ȑ(����(��C���[i*���������AE"��*�L���wl	�q��A� ��Ѵ����(�8�&��|����~{�mM$4��Uv�}���-�n��Ϻ�WX���he�=\�G�eT���3��ދw�%k��s��@��s��l�#*u��OX��3�Z#��1p�1(�n����uyJ%�H���)�Z�w�}x�@��!��U����T=<F�?�������Ɍ)I�p�6��cL)�h&_[���(�����3}�+t�?g1Sᙯ��Er�=��P�#�L��jaU��\m]A)wu�ڔ"O�ܹס2�RP�W>yX�q@m���dW�R�N��[�"\�z�B����)�SPޛ�q��p
}1��"�ձ��W�k�>�ba�s�n����W&�H���Ϩ�Fq7z�mJA��j�IN�z�S��p��a��^E|�Y��\恜ӡ;�y�����&`X`��,yE��`�aT`�oiVw�#(Bu������7��zϠ�!!Xgʌףf�^D�}Z�I����$�ީbP�r0���N��3�K��V� t���} ��|E2(�x���ֶd=+��׃l�C���
E~���+u�3�ͪ�+�~���`b����$n�.B����?���XlxVHYEB    312b     7b0M���) ���:�
6*1q����ˁ���uC��-�%�ыӏX[3V�Om��� ���G.���sI�/x�:N��*�;���sl�K�Q�'��i��֡�55���#�\3l�"�D���ju7*�?�4�h<(�V$�[�82�36����v�Y�άj4�R)�s�I��wU5��Qc��w%���o�ȼH&���S^��Ԛ\��gM��L��i>cOX���Nw��iz�q�lU�UH�H�%�����j�bq������Sq98�x�N��赁C1��m�ojٵ�tedc����|��|K-Y����J�L��MH��%%XzWE���$=_��F�-��ot��A�>���<a )`���kS_�!�
5�;�4�b�^�I��\_�[��5~�N�ﷷ�t�	֒V�}|N��'�G��u�@#�����W�f�?���V��}�}�!JD�l{8x�� ��A8�m��B�h���U�#�z
kg��� o���N%�VX�������)l�b�J�c/SH�&�������`YN���#�.��\�Q&w���,ޢw��v::�?�+5�5$j����ږ��1[��"�`�L(��1�bǋ�]*L@r73���}�ŤCM�"�����>-���� ܓ��p�����Hs���ѵ�XK$�=������1.�PV��'n��;���P�V����T������]c���K�
7p8���^��&H�9X�����EU

�'�Z5���/���m��&)bӷc��%9R�w�h�`��lM�e��	'��6_\?�ZC������|�|�h�T�u ��d9�� ��ă�yP.�`��G�Bl��ұ�����9h¢0wB^ڏ�}��,�u��žT��:ح��������x!����,U۷���>�vG���)��3�d&��,L��t�c��7ZX�¹u�z�V�{�ȌM9)�g�%��!�H1��k�n��\xL���킍�Z�mW�-�}����Ӻ0si���5�X��TV�R"����U����>|Ks�y�>h�8�|�'1��l iߏ��Π��.�@�B�H�}�VM�-�zڎx<��޹�⿼�ߊ�A��y����@��ֽY.?�[�.� ���A�	��H%�h�;Ҳ3G�l�!eW���fU��\��}!
f;��lr��&���Յ\�Y�\�eT���:Z�#]��*��p>�gzl*o<�D(����;�!��Z%~M����ŶW���E�{��(�`T�Lsy��f	v��D��p��%�/ �Σ��(oq#(,�/�����E�3P ��Ngj��f��ߕԫ?7"�K�-\e�q��&5����`�=gL�+��z8E�m�lϹG5�Z�C?.�Ʈ��L�_-���ך7Qo	|�.%_�4�n�o_��#���Q7%��������7�E}���F�'����ڇ�]��Oc�ƚv˒����?`"_�-ˡTR˓?�|�����3���\y���~%��I�
&�$nmp��<�����2r>x��S�S1%0�S|"3�M�u�F�0�7e��!qG����|��xD�sS����.��5�=�1]�R���,
ޜ�@��)9�e�e�b��K}����.�h��
�Lx*Z��,BꈚH)����%S���3/�w�xFv���ghS�����X���A�D'����b�^���4�oE>c�x�;�v�B�T���3�����f�3�|��J>x[s�A����ˡ-ث��d��q�YK��G�z��'��``DM�\si�`�Y�Ƞ��{k2�����h����CN�ȷ���ӡ�H5,_R:��20{�{d���ϲ�):�����kwI���3�^}����XY�us_zĥmV}�p+�~_82 K���k�.'wۗ-u19�' �y���cP��}\��?�\