XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����}���]1�4xŝR�wYݘ������2k�3��������~�;4�lE�j6o�(���6��rӉV�؜�jJ&����erpG\���������3Y��{�KB�'ŷ{|��n�Ɵm�.V����d�������>��,7���4Fgp���S�_�f��D�?w�,"��f�H`B�y��"&Y;���(���QM=�{�^_c�/�׳n4��W�F��v ����%���(h���Z���&b>�=ʪ�D�������-���Rdu%�����i������r������J�r�'������8�Q���D�ם��o�O�i��z�O>Kk�مa?�֮�u�j��n��]q/�]Zb{�M�$��Tgq�W��Hqq���ʀ����uIlҳ������x�Ҍ|aY&�+W�G�I��L�C�q�o�MＸ$�D��(#Ej�YDL�1 �!K���R/ZP�
z�M4h���OL�7fŠ����5�UD��@�X!����U�]��v��d��]`�ҝ�TRWeW@T�&�#[���ϴ���t�kl�'��<����I�f�f��pJ�L~
���U�����`���<m9l�xumkq�Q᪕z_u�����;$�Ǩ9���r��B�B	׽���t�!J�}�"X�?ˌ|�%\.ց�A�K������V��R�a c�N��d�����U�Uz�Caハ�U$�AjV�eyD\S�R�������?zQ��^�^n��M��NJ_����k��XlxVHYEB    41cf     c40o�oⓔ�qxe����c��	��r�dռ� \�������˄�� ��c��ݱ�Y�x�*f�o���E{�c�́�M ^]RR���vԣ�|�T��)����������n��^�0^��~�X|�t�6�����Lˠ��g�����gĎ���~F����� Bkf����i)nR
��w���:T�g�����L������+��*�[Y�@�?HLv���b5T���*�&=�n/�ߋ�8��4&=㱍�����/Ș���}�7���u�u��>�Y�M@0��E�2�sE`	4�:��d���=�t�v��h	�
��ޖo����NH�U6B�d�uRQ�����f=+C�Vs����'�Jm�ވ�߷3)�XXd[�s��	��*� ��p�q��xi���gGbh��TN�Cƍ��Ҫ�c�p�(%S欚�� &�����n` kK�i��6/ ���~�v��{�U�M�fDt}OȨ2zg�ö���������I��}�D���Q�rw��£-�1�
f�4�>���m�Z��
f���p{*Fy"���a�^��YJ�*���luc�m��W�C�rm�~�@���L��n��2h�h�X��8�4ims�,=U�S�NXB�� �좲��gtM�c��~���v"�S��r��7{&�]���
8���Dż$�wa�!)�+��8%&��<1��o�eQ�,��N��������^E/b���ɼ��<�j��5Yl@�?�jbIR��u��Q���1k�c_>��������n����P�h�q��JIQ���������w���-��b_�X��"�I��.�w*d/��c��{�$�h�&%nD��?��R���4�6��Z/��*bRE��Ĵԁ'�A������\W�/�� ��X-��e�'�*�"���R��"Tqf1���+��V%� ����oV��ŚȰ�tJ	n ��/b��-1�+��q�;f�;H䴅��
��̮yzi�ZzV�A�����Rbti�`_�~���~�h|�0]�b+�T6��4*��9|u"�\N\����O�pw����K-�����j�Nu�A,������������#�[���bGA�j�<f���-W5��#�����4���R��8��ԏ����%���0X��'(���=8��/uU(���g@�yPX�F�s�
_)Qt��t_��Q�$�&�y(�d��zf�ͽ?���	�-qh�>)`�>�ѐ��dv�ϯ8��f:h.ׂ1�7u(�,�+�i�[�K�28ټ�K����?�	Eݐ.�
���������,ݏ�=�*�6ĵcdP}UEl|��j��~�ϡ/���n�'��.��8Ly��+������W���O��A�r�V?������W ��랹��*�GD�^W��xpf�z��VAP�P��;���}K���Ǔ-�#!�e��Q�t�燋$��rwBIn�L8�l
#��F��P���E
N.m��h{�ى�=qk�4��?�c�)�`�87����*�x{>�7V��h\6fw?b�ϼ�3��>�X��ȝ7�Qr+�Mg��E<w�F$�y硄�+���2m�'e��T܊z�݄]�j���Ʋ,x�iGl���P�-3�m*�v]R[+Xr���x���3�#���5�d�N�瑦+����K1oU�3�.����(�Lr�e�l��i�����dΫ�]b��K�,�%�&�t�H��<|�)��N��*�j���R�Kd$'�V����f�������ǫpܢK�Ez�
4��Z�K��Ts��P�Ut9!�*��y�̓��b�aXP��#��t@%,��;e�lM�
��'`�%�'��C�*��>k`hT<�ѷ!�=�ּ���"���������>I5k��&�֌63�w�u+p�=vB'y%[L.Tt�M��5���.�����U54F�D�s�]�C��zv��З��jp�������l�+��Ѓ�d[��z΀�P�'�沯���9@��%�����ڗ��ڑ������=�twVi�#�?" �d���U��"��;�O���t�`0@Q�I�ˋ$��ܶCH0�:M7��&μ�"Y�2��G&?F=;&��@\~�����7s�W�Q���Ft�#Sa]��5a=;��T�F�Ă�Dgv�'�1&�w�֕�_e3�3��}��Qq��Խ��%hi���R�Z������Q�VK��qj�j`n|��ҩ2���)�-�S%_����r��|��n�-S�%�O3��A��S~��%�&��r��� �l��_��nQ�C��T�?�����4����״�<�S�q��b���Q�<�ib4J�A�T](?���^j�{-	R)�X9Ǣ��U�c�d��8�!��:H*��B�L�l��>Ӫ�G:L�n������Bʃ���z��{<2��PG��)W}��&�����tL�xz,&�̹v~c�[� #�i���/[.������n������������J^�	�?~?��O]�2\ׯ@,��!�Ě���Jq�z�����m��8�~�����2�2/6�'�D}�
�;���f���^� ]��r�6��#�]|u��)"#�Hʟ�T�7;m���0�;��;�-�W�h���Uʸ�H����׃~T�>�����X�?	��uM1��\�Oى�1�w5���}�6��U��\�a�;�Q���*a[�mHhl�{�aL3�����)i��J3�k�K��d�U�f�,d�c^"�f�7�&�7��[�����@k.I���+C�|'�7"9�,61���i�r!V�gC۶k.4E��wy��̸�Q\<�������Z�SD�
��U^�+Q5�K�RU� PR&��\{�=_z�x�(����K���/�F���:E*X��^�&��4�j ��_`�)Q���=�5'A���q@Ԝt���9R���{�?D���M-q,fܤ�:yh=j#w�"���b����5q�a�c��� ^Ji���(|t��{U,✪s�f���)Ӊ����zWI[�0�]XB��'���b�٭C��Ǽ˻�mJ/n$z�}Ʌ���U���"��p�tW�v�F�s