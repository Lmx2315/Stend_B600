XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��$�r�}.�����SZDr��p}�Դ��m�a}�<���%I��܂��'���+ô��� o��T���s���v�7:*� ���m�����?�\�8`!ņ�`Iסs�H�E,�c���\�*�b:z�T!�<�GH\�3na�9�a\����dk�܋%33Z���S�~G��^(ߋB�	Jp*aoћ��6�x1����G�j8|�	��eS�r���͂])5T���$��X� ��d����.�������7�����v��;��̖�?VH6L��v�e��������q��'7�̪������{��c���P����v�i�}k&�[���z�[E2��]���C6��uD����6�d��G���l�>~��-�K{���x��l$�I�F��DE�`z.� n�թ��zepجJ2_am��5=C��'���#u�˂�g��?Ϫ^4�f�pҘ�E]d�>�@#A�6��"�-�Ch�,�� 5�,��l�Ԡ����U�C`�H
�4Uﰧ}�������oX@��'Iq�=���:�_�=KH��L��"�J �A �w�sG�{)��B����%�v��x>�K��}7R��>�������Ū��a�|����:N��G��5�P(��zͬ�`�Sc�*�5�c�����O�C~�'f��
����WZ#�����˚��C#��)��ݘ��4��L���*��g�fa���G�Vy�p'���2U4R<:�+��ؚXlxVHYEB     6c5     300��ua��̷��B�p�t[�#��H���v�?cw/sy��z&(����˯��0�����,�6ŞJa����{9�d4�^�;��udmN)����!�_�4Fغf�	�z|V/a��!u�<(�a�1��|Ɖ��s�3*`Wϴl��6���h����FcMLA�$�#�"4�5��I�b��G��������`���.eh�A��Tk�j_�0��xf������͏�vi�:�4�*p�EJ{1�q�ͩ��
���s���z������\nR�2��E��i����? 4C(rKz�ҹ���f�wN��C�����-��6B�U�����s�oB�4$���o#�&	4���r�mg�4�@=7=P>3?Q�����2Ki1j�l9��u���������S�Y�@��Y
M!��ry��)�%P����A/#�*F���R*Mz���ӡvvЭL��<L��D���Nn�~$�2�2�ms���)�9Z���(u����G�Ooq�E�w�)�%�$����aU�J��v�
Jb{�C���iZy�8�|)s�;ᗝ�e��t�tc�A�p�9
�Ibp�W�H��~!)'{�n�2IM���w���Cb$��H�7��;�NM존@qJbGVj��^'u/K� ��ͯ���x�OΖ�oU���:r�,T���K������P�o�9�N1T��EW;D����KP�(��� ;���.��xWN'ϻ|pjs*�Lga�@P���jfn��7�f>t�ťp��L\_H