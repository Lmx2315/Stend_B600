XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���/3�K��7j���H�=�/�������������o��js�P'���c��ewC�߅A"������LL#��و�p¦Qw�K����bÑ͆	v�����;)ћ��=b�d��F�Ot��k>ڒt�&ۺc{%lLO8�vp��� [�z�y����/mX�� W;�%�q�&o�EΕ�l�
������I3����ۓ��7Y H����,����o�CJ��+Tq�>�f�{�O|;��Z�b-8���KPD����Τ'�'���?ee��uo<��|D�lw�����u��RR��9��u	��[�h4De�����"��e6��+�'�	�����/�>�m�:�Vf9���*�l�1?[�^GL�L�v�ܠ�N�s���VػT�3�q4��/�mO�YИ�}A�uYs�.Cޗ���;�|t_���^�4M2���~\ֵܿ���V\�����]L�F�ld) �rXG����[�qo�_ʊ|�f#����<>�W#���gx-::K�'�kX���I<��	��,���<8Y�s�c�GSP/݋V��bo"�9�b���������],�Y���?�	 �BM���IȌэ>
�'��~G)���b~o}��,���'s�0��t�G�������i�Q���%��-oz�bS�a�Sl�AM�ڷIŴ��"_�p-�<I ��F�G}�?�F����&���PYO�,�<�׎��k�+�����P���W*/�XlxVHYEB    1901     450lă�u�-�����/V�4H5���+�u'6+_/�Nz���+�^���R��������J2Q�W�sM̤?mD�T�����,1�f3�d�j����Nz� �l���B3�<o�O��[ts�u�1�d_B��Y���\9��T#xX��8_��ߥ ;Π�3�0DW�[�X%A9�tO�F�X:/�܄'s<��g���7"*��H�(�e���m�PVk�����fli~"8T$>��/�mtE�
�6o�ygy�7_�s�wkW)>�% R�>�qd���8ҍd����"[����=�mۺ��5�Y7t�1�,���s�`�\�:��3�t��i	7���7;D���-��5	��/�>��Z�\)�V_o`XDԂ�Z{s�;Ϊ�r^�g��	'�8�p���h�{G���c���68���b��u�[F��X��	�%2	�.>{�WG��w���<>�9=窼�Rj��3h%����6#|L���H�<*�z�V��-ߒ?aV��ƶ��'��l��LJ��<��7��ysɺ&�%E���m�6��)X׸�.}9���5�{�':ɖ8��|�3j���+9��^&}��m�;N�!U�By�w�i��{�)�<;����N�'*'�X��I�v����5e�sn6���s�xF�]��cJ���v6�
/�L���$��s��f��~
�w�%��|n����؁�}�x����:V��r���QfuP,�wL�y��~wzb��Of+��ʡ�wL+P(ǴU��њ_�~�ya2S��d��р�P����5�D�耟OX���|��	�*�+Fl��(�~$F�j��\�o�\�C��1�EСB��p��$r�����I����:��jT'H���Y4�"/����<@�h��jDНmR(��f��;}��л�M���"=���f�o�&}����ʚ���@B�i���i�P~����7B�rQ�֬��ID�X'Fr��AJcf5��3`�PZ�Ӫ"�>�ޯ:��Փ~?%��Q��LM�$�! =eI�[ �r���:��5��8/��]ΌOJ^b7�*;���Ԍ-+�P���+3�A�m��W��ٮK��e+*