XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����q1-��KVն�C�s�R���ԃt`-�M�Kd�I܍����6 ��ҡ
^4a)�ML57��hmȸc��OV�r3bQ�{���@�)��=מ�	A�Z��������{6��t ��<�1�0<����锗�oV5�kS�r,{V��}�K�W|����4���j_��Pgns�#�氕b��4��� 0�_�M����AO�=:�<��Njv�B�6*5��9:#��.}��`l��F�@�
T/��X����5����;�A�sZs�FU�'l�M�B�) ��nJ5�����u�7�T�u�̬�I����Y"�a�r7�o[I�o=����w��|��FTc�	��Z����m�E,7�ƚ���!��Ԫۭᝠ!4<�j�]}���8�ۆ��=h�^��K���	~w�D����,"�~3IU,�o �A���n�8Gj@ �.܏�˴��R�����ޚ�n@/4pʘ�㊳ڢ5�/������z��Ҋؗ�����)ֳZ/?�f{i�%�?L�������y��h F81lH` �4�e��V�WƀUĲT0���l�y���]��@�v/��wV�7
�x��X�1ѫ1��øt�W�/o�����S�t�h�v+&��
���K����1�f�IV��"'��u!dK���GTOD?S��F9�-�_,�[��x�£��g�.����=���@9�`~�$ü��d-���d���ϐP�;�j��󸕑Ǫ{�|[�R;�7����3v�YXlxVHYEB    3a1b     d4041��8Hyß> dՌص �5wp}D�?��$�Xa����B,��چ0�I�c*�~� v}��B��(���>=��M�;��V�qe��"O��j�)-���,��㥪����G5`5/ ��&��?x#HP���<�����)��$e����v��]V8��Ic�
�Ax��%�����I�S�L#y $��R��+�%�)6C��>�M�ȝ_/rIeK�=��/@y��A����Q��#<�v��yj~��z꩷f._����x��\�E<�v1�D��t(�d�cs��Z�6	Q[P�����v�PH��Y���r�|ǵd�Խ/^\����dj/5�s7��
���r>�����s����)"ŰDS��=pt����[��@����nr�zIc!�/�X]����#���߲����%ڈ��Hl�)�G��a����]eā��Df� �6��L֯�:I�|�ac�Đ��-<��x��|:c�!F�3���@bLg��M)��ot�d�p��i���8_l�$�t��Oi��3�����{0�I'��%$��Z�m�����P���<��T�-���L�ɖ��)�]� �)���\��%��kw]Fp�fa�V�1�CH�k��3D�$BA��T�Ϻ��{M�.%�tf-��  �������0��NaKL�����;Et��㽣k0�	.����8��$��/<�>=�Q�N*��P�.u� ����*�ۖ}�wL���:d�=D�q�����~���v��>m^b|Jt�<p��}�!>"G����J��yGG��R�:�J�6�S�^:O1�f��Z�T���v�d�_~/�� �C���Û�����\����ɝ�ⱙ�ծ��e5{�
�+<d�n��T~xYȑ��/��'%�fJ��*�i�R�Zhc� n���E�p��]
��ۃ�1?��9�C�p��#�o$�s�������
��m�6��筝�;�'��0F�����m��8Nur6�2n�u�e�k�	
PK���'Y?f�ե���jy��;�ͽBۛ�]�(%��)�5BT�.����q���{zS�>��>~ˑ5m�JW�R��89z��^q��m��N33*�ȴ��%E��(I�Oq����*-W�`Y7׮�����p/iQ8�|
�V^�Y�~�d؞g�H��{����<�����'J?����,�ퟪ<��k�B��ݭ�jzF6�|�Vڪa��2d�����1=씄��ȴ��T�LP�����mg���f�n@��r��(��p/�H�Ќ�)	X���4U�X`�����kO���@(���8F��c�f1��5�%#8�i�ì���cA���xa�;<������<p7�	}~=I9a�1c ����Mna�9
�i8�P��5ߧ��2���!��nD�o��Ϸ�f���'����k�'<T$���F{.p�Q�ˍyx�Gl�<���u������S41�_[}?�-�l̣�Zܑ7���A���vę��-fH�]�*� "-=_��T���ş�q����N 	]ʑȗs7�H���M2��G\�\X��I�*��*�ˮ�#��}���Rz/\��soxS���mW�d5���/5�ޚ0b�U��Y����4h2��k`�T��Y	���d:HaKwor�j��Vp�XW�B����^�<=yNc�5�.�X�[��Y���s�bg��TZ�]Y
)��Ѓ��y��ŋ!Y��7�r��Ѳ��kd�C/u����<P~	��U�t�Nh� ��l�֫�a���7W��@,��^���1�u�������I�� ���̓M�x@���ѬY���m<����oi C�u��r1����P<�IL�=�3����e�#6I����_Ke �B����n�'�M� �	�7�[-���Ă����a7�T`�� >ݑB�
���s�qEB�e8\�'�l��V�8da]כ�]�TK ��{	�+n;�{R��%��p��{w�&�l����K;6�S	@����e\Q&߱g��SY�7��X���6�l�Lo��M��.8K 	y*����ߒ!�=oBQ�i�ř���y�ơ9��0=�19
'+����V�q�mݑf�!'[%�=Id�[ꚔZ�PzCAc��h�i���3���U)��C�K���ԓVY�Aقh��9c�mW8�j_?˃8̽Q@�"O�Ӵ��
�d.:�BT��I��5t#��$�xDuۜ0aIB�z�m훥2��v����(��3����:�X2>�����6��8�DWlAP�+� ����Ekܛ�Xxuzs�]�0��3��AQ��ͫ2;�E>[�{0�Ù��n�<O?v��4iA��OJ����+�;F��	ff�}̺�o�!k ��FfбPu�*�����A����P�3p�l)D�W�B�d�XNv������  J�>�H)�Wʓ1|�	��ݻ��\�L(�c$dHR��1Wv	�o���y!��M�/��N�Ώ�ˢMp��J]�m�ڋ�d���1:�)�w�)�wduFT����ܾ;]C
�8}'�N�s�H��:ү< � ���>`<�xc�lшz��~Χ�"=�ZՖm���e"���	rQ(ZU�0{��k��3�>q�]1�%��� ^�Qi�
�Ȕ�����&�Qu036m���A��h���ngBW��Q����w����?ʯK=�h�LT�k�ئ.$��l�Q�~�D�o]��m�V㓨!S(��4_���s#�V�f���D�foV�q�-;"�����z�Er�z6��9�k�gGD��%h-+�ɻ{UߴcK�Z���H�+�>M�0��G3{��j�4��	_�$������^�R��|�j�g��-���"�y�j,�`��0r�"��S��E�C�.��gb_d���%���)�-w��j�ǝ��+J�}�����?V���C��P����Z^%�*�U:�@T�o�T�,y�������ZF(׷|�^������c�&8�����;ڗ���Ҿ.�f+�#h�(*�dzg�_x�QRZ�{�X*-D�J&�X�FП1�6�
i�{:�|�z�f"�q��F��H�o�߮(��2Qb�h�L�\�<�\��\@��Pj*�#�Y	NנG,�%]��{ӄ{}qN�(��r4=��\d�|�_5�R�#[�=�(���G�X�R��q��}���Zvn��������vl�f���2*	�ѷ?��:��t����di���4�y�����%_^����{̱�d����$��^m��:)l��fJ�'.���?��Y�ƨ
55��`����'_<�
��L_ywSu���|�NnR(��!f��A��gEr:)/�vQ.����G r��9�7*�O�