XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����%� ��2�T�<�&
n�-�z#ݥ�h�@�,#)y1֘X6�j�uY!sk���:�/,u9S��cJ���s��%]QKMJ�8=8�O�*�qwB�!���7�$���̸뎇<�����G�ʊB�P�H|�<5Һ�fҦBeJ�������t��� ���L�&4��gO7�6���D�Ôg�RRgn#�x1/L��f�H@��	v{���#�6�B�g!$�s�t��C���f�*������m%B�����rhK_�K��A�RB-��Y�V��Pq�bsn�B+�$�� "���o Ú�'��ou��Ӝ#��S�*a��^_|�UN��������Q� ��/�,F9ş�/��-`��w�pɔ�U ���.�]�Jg_P�ZƪF��mcsc��/Z��jb���YW`/��2g���O�M��o�Ɨr��̹���u��d��Ò�0�$�(.�{lZ�CS���Wc
訾��9%F��Neأdg(ig�~ ���Ȱ��
�S���9n:��-ϸ��!	0���}�6���zc��*u)�H�|lr79-�4�W�v�S =J#q��]@OY�{��Ł�lhRU�n5���TRm4����,M4�~zF�����E���&�0�l��b@,���j;$2v���K]��{�fYf�ұV�jtW�E�������/Wc����)�����@�rW�ufO�(����R���ʛvB��`ɚE>�>_�e?�5���P��#?�8ӈ&���q��=R��0�I!;}bXlxVHYEB    1578     5a04 �:r���b;�0f;�UȨ��ҋC���ۣ�s%���T�Za!�e<X��,�@h��v]g��h�7��6��[z4�:���U8
�f[N��'�<?;>FDU�2?�`͵N�N�+\��M��_��5��?��p�ܲ�-���ㅡ���+���J�:����L�Yy�yؔ�7�':�Yo�B!Q�MN��N�[{�)�b����W0a.�n.��t��n�M�F`��@UFr��.i�ʡe	U-��]���;���?����ɞ 6�D��XN�|�I6�k��]_��~_��
�,��p25'�w ���CG$�h$�ʈ��赓X��C��ڡ��u�[��'�c�����ێB�|N��9�=�,�qB�(x������z�+
u\��I(�P��.��� ����M\]$)�lT?���O�~�{h_��fk%�!!��ʹT5�'������G]���u|�s?l��7�,� F�J�S�ޱ�(L��`-kT�λ�a*��S�wձK�
�Y���1~�C�mZc�n��%���z�Jx�N_�h�ڄ&0,�{�Xl�b�b(�c��}�Y#�W΂͍��$D�ય�/��f���ƼkZ��6HB���s<J2�?�
7�ߪ�6�&(��ǿ��l�͗^��90�fw�v�~��ȓ����ޑѹ�]~��P�	�>0��ӆ�~����U~�"C��=�E'!���O�d����!N��`-��i�(LD����;�οd�2���^�-"�V"&�6�Q�=:�!�K3�	MǶ��p:���W�K�w���F���B���v(���X�����f���$,2m�_���%+�9@�:�f�Q]��~��IT�?�0��WN1��=i�2��IL�,�2,W�)'ha��M(-�y�@��W�a���o����)�-D�� Bo�<��l`f���{���hQ'� ��s��3@$�J/#�#�>����=7nG�8���Q��LC��� ՚�������i>�r��d4��A�t����BC�����u6|��.v+kRA�o��{������\�g(y���w#��Β�k��C�/�����̦6Fs(��@p��73���*�1�X y[���\��Ƚ�.�4VGDϥi�(`��x.۩�Ke#v�-�J������=t.�k��m�'����|O^�Պ�y��_�(-����*Fr]"�6�1P�#B+@nN�V������Y�$�'r��<�<30��ھ��V�Q)r��?z���0IneF�BU'������ˣ2��`9��ᥡ<��\/�4Ƭ�3�i���5��K�Z��ЍeZH������)CYx�|Y�M���d���'�7Fs�`�g�9�m��le̵׌U��'�,�7��p��zE�LG=ۃ(��͉:��F����<�f,�I������2G�