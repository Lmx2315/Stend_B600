XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���zz$�J�4Z2mh$��>�B��da��]]q�I� 4ry��"͎���}�Q6���6#�/�+A*c.����r`���x�f��l/)D
��	+��rD�=�B�4X}��Ģ�𛿚u �[�e�џ��,���՚'@��=��G��J��-eO�7�2�9��
��mw����(���Y�@4���\��U�/�5�57�+[c_�B�E袾W\����D]Wr�&�$�-�(�mJlӀ���?�%0H�6�bM�����%"4����f�,�]e
m�NI�a!���w=�L����Lo}B�!O3�c�MŶS<4L�w�t#�c"�j6�\b����rO�3���[y��>�3��|+�a.N5�1#u{�x8[OI�-Ҁt�|��Sm]d|�����tD��
�7u;]f(J\-MoҨ��(�=�7�q�J!�]�]Y�ePPqŏ��+$��H��a^%�؛ȋ+�{{�v��&U�2�.���9�����yz!���lO8���׻�"�����vv~ �CQ�'n�1�S�����e��N�c��+w��]���T��n�RF=��<_:��!Zۃ���ŴehV��3�l蓪��ø
�3�X5sӶb� d��Q�,�J���90)�15E��u��h��F>3�p���V�D��Ⱦ[+�����q	�˾�G�z�J�
���܌��sJl s��� Hk��[b3�'�n� |KK��V,�/�(�V�~��p���]�n֬��ߓQ�D��LP�GM/�GiXlxVHYEB    3246     990t5R�
/�Zp�t�L�e#�V�3��=%s�Ȭ������SzT��)���� :�������?���Zl�,h ��c�Hf`��r�S��p�,9SX9E5W9^�K]t���`@_I
U�W"���Wz�y�B�Yy�H��dq!y^y����]!E/� ե��o�$�uLu�3[��s�ڃ���`��F�^[?���P��R��Qu�8���B�����{ +�Kk�oO�F�!e����E��RW����n�3�����Ŏ{d	]o�)L��F�^"��^��.~i8�F@޷��Z�峯�o]b���t�J˒*D
X�J�$Ͼ�o�(�ڼ�#e���>Ӌk�~҇��t0�� �����G8�͗���ve�X\ꦚ��R�O�urM/qd`�C!o?&�|[���`�Vu��\e��{vʫ#�������3'��y����vVTc�B����W�B�po�S YW��p�#u�!��e�/��<n|�&�c-�j���kA��Tt�)ȴ�~�J8�qѲ��4�x�'�fi\��ZQ�V |?Cv����W�O]��t?F�;q������S�[w	��|D��3�x�򧕄�X�uUBV&i�bA%�{�]�*�r1��݇���������Ev���f�]^�Hw�C&��%��5^aFLQ=�}��^kL���Esԏ`��
�����]�@A'�A�@bŘ�"�}'�K���8ڃHG�)A~n�%�N]�,���cz���x��a�ը>��y���=d�"��E�����J!��4�������U$�^}Z����?���&m\��
x5��ܻ;��Ә�Ǯ��P�6$���z�3�p*Z#x�?��S�e�Ƣ~���(ɐ����Ỽ�g_��/t�$�3�����ezU�48����Nԝ����6<$��uU�s0!]�,���q��C�uG��V����b�R�/������K��'�-��^�T�WCE����-���G�A5#%T7 ��� #�(P���rĝ�[�Te�6��#�O�_�	�f�B;w�X'AM0�z� �Y� ��bQؤ��\�
	z^o�0Ǹ� �e � |�xLc�J�d��(T%Ynb,2���C�r����5m���������bwmr�ZV���ݙ�'�����==]=I31O� N�����S����k�{7�K�y�c�fD�����u��2�I�0]��< Lf�����nH�dW�Mm���z����w)�Z��^�$஭��������m�>\��
Ā]YJC�+��W���x�S^�ЏH�H�9����a��#�r��H|���H.dד�S\�y��![���Y�K�(�Y'�Tx��mtg�RV�K�vj�ޏ�w�C|t���ƷOU��᳴�OE*#~��B�S����)d�Q�=9�؅��.8�,�A��Rk��$�_���Uy���D�����,͸^���`u͗ܵP&hx��́���@v�-���KU����$�$���g�7�>e���pn��2��MϜ&�w8ws�N��P����_h5���A��H�(w6V|��`��q����M���}޻o�]����F�
�u��V��~?�ġ��	�yf ���B�I�ԧ�=1�O�l��n)I����qݕzlm��:�tc�J2�@hH�ը���2Ф7S�ͱB�0�����E2GZ���x�F�o-F^`���4J�.df�����+��I/F�;��.��1�Cq�h���#��5��<7�!��%��F۝�%)��J��֨�?@��5��2�֕CQ_[	]DqT�]�b��Zp>�1��97-딱�{q<b�n���.$�CL~�/Ẇ��\n6CNWN���ueH;=L)7��XU�n5�2z#�<�֪&�ٵI��y���K8	`D��0/,u.���[�r��[Q|��O�}�tM���N��%��f�F׉�濊�,�k~��Aq,T����V�Od��$�Kt�xĞa�9��2 �X�XvS蕕��.�)�s���L�6�r#F�m��1�,�]E@�)�i�HW�v��zTC'8���XW�����Ԉ��	�8o��z�Z�q3�ȾFVI#��ITbj̤�J������P
D�/a�z�'�ֹ��P����d��,��f�)k{�K5}j�z�d:��(a���j�J�&�a1_S)���.>TC�C��5ƽ�s�w����E��d]qP����i.�Z�-x|-�4�Y��-��I�B@��-�r������pf�BZn�֞C���ʽ��_����.�Su2�A�>L�����m��w�*n�c	�"�'ہ��A�s[t�fS��R "D�
�_�����L����d���;'j�R؇Oσ߫	�mD�c^M�oβ�2�M�^�c�"o˹@�p9$�v