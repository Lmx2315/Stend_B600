XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ؗ:�;��m%�S��w�x�+��Y�[k�\M��qp�λ�����}R&m���������-{�C'��cTm�ȪK���Vs ����o��ѐ�uK���ǂ���3��p`����MH����p��$��NO�9�wV|����Mv�k�B�����1�� T��C,{Q���(?��?T��0�
A
�ɣ�4� �!n1]����87���
 h,�A����󝑶ɸ	GH�vL�8���p�~Nn�Z�y�.=��.�"{ŤH��.���r�g�P	�(V��}a[W�b#~$_K����8��"�ɣc ߲j9�SZȿqH�hc<����u���JX(Cv�4F�ލ���u�_#���s��V�Np�ll�#pC=u�O�r�T�+�|�0��"���ۛL��br~J��c���B �kJ�GU�5��;�]Z%��&U8>��V��Ŝ�v麯��Y��� �!��l)G ;���F8s(���8�>���ؚ��Ke���9�N^)rc.7;T���K}�<���{�Yf�Usw�}#<�lj �f׺���`�ZN�	�����q�%�����V�~�[��w�������7kO��[�2n%y�����I+@ DS�K�sĄk|mxZP,Y���[���Z(�I�^�`�0�
��m����\��y�xu7�0��"|
��n�<��iF�\��Bu38zj:��Ϗ���dnn���u�{��v����'[S�D�dXlxVHYEB    1046     4a0���)�z�&���T��*|p_������2b[�����>(ۍ _J+��,3��|������uх��߇Ӓ��Gv��F����o���0��0&l/�}�p:u8NQP6�;�����	�І�юu�Ȓ�=�B}�a�q��<Jv4�$���Lnɟa�̘�,(V��#W2Sذ:�V�`6�m<���M]_��=)E��T����XEĸHy7T��T�ذV�����\�5	��Q���c��x�"�� ^�$|��'ﲕ�Oc��a�t��J�����9_P�^���*Ϝm`����1&�#��p%%�k�����&9�H�>��B|�����.u,9�5����{���H���:n�bA6 G-����gcc��;>�J
Y�(���7��©hb�}��+RY��v���R�C�1��|]�Pn�]�đ�y������x�3���/���)Z��s��X(��٪�M�l��{Z�H0�2���<��zJ�"����6.��P�V�^b-=�ٜ�
1�@Kܥ��U'i�2�W�ɨN����I�Ej"��04�5�� 5۷�C��SC,�����'>��=�p��1�:I>V���k�^u�Lz(�άҿ�iK~6�M�+���J'�;D�8>��4� 욏9�c���Q-��|SIX$��z\�h̚^���5]NuR|�V����D�"W���6���a3� ��*ɵ��Ӓ�:EW哛�{;h���z3�r �"�qSz�1FP�T[R(�K����6Y[�zc�"B{E6�D����ª�IVD��)7J���*�r��&npcz��=Z}�gB�?d6�2�l1�/s�g���.��0Z�s�j]��z9�J(�쏢9�}��/�)��H�����L�b�_PĠ��Ci\�e���*��V�A�f�;��a�8�h~��	K�/����Ol�-*��z�(�ɧ�K���qy�4w;�ߜ:j%�XGɠ+"��	�m��yN&@UR ���2�7ӊn�F���Lp�'�*���Jλ�v�ö���5�Y�e���5
vοj�D���s3�x=T�z�!�[�&oH�a�[-XF�c�E=����D��^�}xH�B��(�2?j��0۷A�i��"�Y��O�����'U��-@􆷴�Kf�ɠ�}uI�>��