XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���q�3�ڊV��aġG�z=T��.��4�ڍ����Q�
?�����U�@�?A"�1ͤ�)�SA�z�� 	e5�hx"�j̍G��&�����j���Эۭ�� ���uR�\K��Ø�_WX��u[0�U�w����L�)t����ȋy#�Ԫ%�
��B����>�4}3�l�7(."��+�qY��܄_vs���9=n�e?�Oe�Zgz�Kxɶ�ڜ�]B�sq��� �'1�!�Qޚ<x�C�шR�m�f��MP��9�i���NcDk�$��#=K�G/�!�ƺ�{G^>���"D�/b�.���n��/{\�o�Y$&g$��ֈǌ.�]pl9��p���:Jx�Z!�B�z��[��n#���)�'��d����ȿ�Ͷnt[����'�כ�.W���q���S���9k����J��Cэp��|j?Q�dk�.,Iz�1�����.�~|)��d��Y�,�J������{��~�D^���*7V�0�U���o3�Y!L�b���j���w� &흎���q�3~с���(gyx��V�`'����q����^�2jp]�K�:�W��+��L!�P��1��q�.�ε�OtbB͜i�Ѿ��'���Q��T���`��o7B�n�nj�hDN..0��sPj	<`�-6�&�!B�SB�#!�R>���4:ؿ��AJ
!��?3 �V�B�r����!y����{��'��.@���XlxVHYEB    7e17     de0�vXOE�?�&��j��X�!p��<>67�ȱcv��=�8��2�0w��P�[q��=�"a/��?L\��B�u�ҧG��U��ڕ��[�@4(-��!��"s�rF�>�a$5)E�c���͊�E!������H���A,7��2o�+�w����_q��Y�㾮�D���q��=��V�+�E��Ey�['�Yʊ�V9ω����C�q�Yl�k��{��Z�y���ݤ���R���ik(רX7�mTV�W:,����T?{!ɖ��#f(4a`"�֘�F���n3�|0
~I���/]XY =��`��j>���O�3_?�0�	T�j����6wpJ������n��u�U�o�1h��@𳣢թ�g�,A\cqH��b55`L���G��Bb����k�����'�篺BM���i\gr�XBh�ǧ%�h���R���)�F�h@�"��J�_玲����J�͞5}��a����e����?ƾ�I��7�R��f(e�I�`���5�n�[j����x륫��'R�M�
E�j�]Z��OM|^WKЀ`=O��:�� z3� ��}��s�|"7Y���+�Õ���t�4��������}�5,���|AZu���x*/�k��IB�A��.F7֞o���.)E��x3(�q�(}k�SB[lBw���B&�8���_�_���v�W��~���Kv{��"v�6V$z� ����Y����W���R����[찡%��\:3žU�i����R��~�0AjZx�( �C�g��e!7�����#fe'&$��nǟn\��̂zK�����>��
3g7/\��!�[y��ΛL�l��0L�̟ �kY�R*5 ��6\�R �|1(Ak����no�.[��x�CNol�&�47:���	N1t���2�lB�"�KN]/�U�P+QP�';z.�8�� ���������Uz�A����z�u�e��0��)PM2S�����8�����G�Ӡ�jb�5�q1��Q#�2�i�x���{�%�Ε�%�#��G\K���m��4e$@�����e���O{P"�Sefj@F�E*P�"
���<Ja
(����E'0J�������̼��p�VD�����@k�]��^��`:�wB�f�A�x,9�N}�	��ٝL�>2�&%@ � |t�%B�}.pz���ǐ�Q��Ϗytf����u�X�y�z���	I;5�,����H����R�N�|�:�:9T!(�1��)�#��4o�j(����f�vi+�"����r���i����)|�M��Di�%��q�⛙�Zn�i��lK�>�S�)�l���9��b���Nѣ�)q�b�C]Fs>j&�D�5}8�kN���p@�
�e�X��6!�T�r�=|�0�T��3�v۩���hP����`��0�b�+.u�k���~O[�w�U0�,���ˢ�&�1V��|����謧��y��^�HE�1��턋�R��0�x���I�������Z*!��Y�� �4��x���F�~���<��S�R��ǅ��w�d�O/��|�&��q�r���S!��a~y;�k��@ʽ��q~����\'�j����[����K �;��a� \3]#���V�ӵQ~I���g:qW1�}I��p�(�`��*v`��b��N{��Ǳi[��lQ�T�u�y>���.�W��H��h��Z�ȉ�8JB���+#��ˎ�Q��#A���@3�;�'&�SO�]����Ė#�_^���tT�;�]����]���.�O����ӂӢ��2WY#�,�爍����{��w6�j�4��zqPH���i#�X����<���&�HsV�)}r�=��[����Ro�zH��s�+ϩ�,��;���Jݛ2���G��h��aSm��Ň�U��~��nu�X��
�J�}�k�V�dꖭh(�Rb�6±D��ہ���ق����L��3�`F�9*b��E ���T�Ê:��0�Ws:�]y����E2�V;���;s��7
 �k�
�sQL�1��\g �X�����4(Om\R-�a���ӳ~�l\�#.�٫�,S�Ka�� ;�3�\	e��ȅ%Jd">h�������t�di����㿁��O�w�ơ�Cw��y�p����t�Xw���I�PJ?ߙIUv�c2���R��ލ�s����?=E�
�
��!����`՗�
3P�y�A�%?� �s,o�G>Q��=s���d�4n\F�珲���_�V�6�}�ط>{���]?�N?��7>W�Ϥ����HK�'Re�iӕ|%��l��9�*Qt-�f$�E����N����&�0kv�$4:���<���}Û+�,�#N\x�?b��1�#��0���1&��6��߶O�Nķt�5�?��s����w������ꗦ�GF���+F{M����)�ϻ��>}G���Q"`�hj�>�.�"8�oz��ěp����(�����6��/U�����..��U��</W��{Ǝsi��Łn!�&�&� �4�U�}����؜=�	�z&���5�P_�����e�ٌð��:��-���_�Qۭ�����kp�&Ϩn��Z�О�#�?�R�@Jۥ��ǣ�.�4Q	��z��B���_�Z-5��x�HiB'�ഫ�Z���q���
6	��Ƶrx>=�2�S�'U�vO]� gm��G�=u�_���Ù��0ܨ��"Ͱ�ǚի*��+W���k$lS���!�:��Xq{�� �}P��Z��4�BPɮ˭&�3qG�wQ�u��p�01����e�6��eʝ��N����e�/;+H��f���d��{�U�p)��x����6g�zX��*����~��Ɖ�����Y��q$o�Ą����4|Q�#�<���cu� ��A�k ��冺s:;ξX��N�F�U��x�jP!ldUA�C�������o@7���(��R�G��p��}���/�d�깜Vػ+�l�a?��J�bD������ؾ�:��ZT����4&���y��X{���ʬ��7��O`w��v�`���*8�dc��l�2'5���[yG�>��~U�)������V43Y�:�h^o���/w[$#��|����� �#��r:Bx��z�i���~��2���Md�mv�0I�Z燶UQprԴt�0�c����,���p�\i��@	���p�
����o���@W���9n̏�"3�\�Av	�n��u��߽���Z�J���ޠXk?�Q> �]b��56D��{��
Ģ���p*9��^_��^x�7���3����L�{ C�S����;iP��;\љ@A�S�eȫ��Ш��ͱ!�<W�V�F����,��kyX�AC����534����^9 ��S�b՜p=~Σ�+���wJ��[	�(R�BV���|8�u��<���l�I�mڑ�a�u�.Kiv��ݞ��`�zs;)>��`)��=��쫖��0�