XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����K�7�M�t9#��۩I�H~�J짉�ʇbZ'j����M���&���e�?��_.&���k +
'�,	N�{��A�;}����#�����6�Bc��XC_�
x\�.���Ҫ[3ulq����tmZ�ڟ2R@�>�oB�eh'���ފ���g��Q��9wWol
Y�"�%MM)�ݓ�z��*����ʏS�1�JL�Tf4�`���B�+�T�y��0���%���J�k�]���.|���۴(Bk͂@g����?��>H~�a�l��U�ԟ�4�i�������1GetD�!7:�H�m�N�/�	�u���^HE����mc�(�Z?�m�s����J�ȿ��<���	�"����}�|�ڷ���� �D��΂/�AB|�%k{2 )�O��`H�uk�?�5�9|2���}F��Ն�7�~��c������V0���u��q�c��&?����jV��a�f�> �N��"��E��h?ֹ���@�J������/i>џ��}��o��茫��?��38����P~�.1j�F�q����P����2h��Q8J�60Ȗ�ﰔ�gՠі[B�u �(&���p�&�He�@�m^�.}���:�">��OQW�C=��S�>�G��8�6�i�`�9��?�.���R�L��g��P��;9�ߖ7�K�.~i3���t�` � �WQ�1�'u�V���^�DM��0��tPb�:l����}��eW������bzpd���95O�\�=�V}XlxVHYEB    1041     4a0Nqs��������*Qkf.�?��1���zWѢo���_�;k���˶ >	���s��!�9�7 �Ȫi0�=�9-G��� �OB�
��A
����#cN�ST-y�w�c_��YD�
{?�OS/��K����ͬ%��jb�S�Mu.�+����~jO{=�Rd�9��0�D
u+h��_�!!�G(p��u����s���� w��ԙQX�xG���K6L���݋�c��J��&w?�Wk���ٌ�1�7�n�i��+��L�T��Pƪ���B?��Pa�ْ��V(��2�|S��z�A�O�{�g�sHK���v^Z�uVqr��Dh՜$�u̺`���|�}`��ո�����&d�@�gHk'k9p ����T٬������S?ܝ�����o̜���3PR0=�'��o��>��'�:�h���(�f[t9Q�{~�uķ�w��f�"�u�Ҥ�'�Q�|��B��2+�����b����r�[�s��=Er~%ߙ�|�B�Zbg���}���c�G���h��T�	��M6�}\(�<'���ֽ��ND�]Z/���I�3SP�����r�H�n��}({�Pc2~���`�a��8�+��I�����W�m��I�A�q�7��{īg�>���:�@ml�?4�1~`4�"$]~��[���QO:(����sk�Y�Dω�U3H[n	�}T�%/�wj5�_G��j�$���H�$�'�bN�ArCB�;��2��M^d����K�
m�-�r�~�[	!+���h��_~/��b�r�P'o�ך������3����o3J\���Հ��㼜Xz^���D_ЄmF�y)]��Ь�(Zr\]�$^/;}vn�@t����
ɮ&�$^� �r��=k_QrH,p֡9S����]4GM)hᑛߠ�eg�̤ۭ�dD�@�G9��ks�k�<A(�9��4��Ꟍ'�g���I�^�1���d`��Q7+l�h�pKw'��;3�s8}e��[��"x4���4l�A��Kt���aZ�p|�h�ħZ�de�yخ��_cO�Co���3�!�0�7�<�����{����9Q40���s���] �Zz�L���$V��h���|�>t\��抜�6���$ X�?�gL�]`bK��ۤMn�.�6�\�ђ