XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��G�*��q��V�tO2�˽N
���S�z�L�"��rCvm�`���lQ/�$�����}��p���Ū��1�R����4�����1U2������%��^1/��m�$�
���&.Ө�'�\��*�+�:�7�lf����E�됯�3j��&X��QV_��h/�N>��AƒQ�KWj�\���M��d2����s��O��PKޛy2�a����APՀ��O�d��X�Ԩ�Q�O�6*9=�¸6W܅P�
Ov���
������~��#��3�j
�{�ɱ�<6�ߨ��@���'�����q����K&
�h�"Q7X;Pc�l�)�H�hm�����̲�ɾ(���oj���?> �aי>/��5f[Ŷ.�����
o��ٳ�P{�y��М�	%qO�h7�B����4�!��	��$�C�p$��ɨ��AZ��a.M��2��X������w1Xc~�����14�/Q�C�b�	e�
2�Ѱ&�Y�$����uX�g�Wp�N���?n�s.��+>����c-{'�[*80I��ف��=(�5����u���6�2��4�����g�w?���$�@x�T�:Z�my���J����FM�|S��XR>�%%ި'� $�>�:���@��Ό{M���qB�"��앵9���-OҾn2���"��H����%лIu*��h O�.�2�[_�9٫G�I�ZgFß�/��R�8�ǇU���Y)�\� �����׎I���ɊXlxVHYEB     748     310����YF��j���ۉ�c6�Y1�%Nڞ⟈��h/ѫ��?kӐꚮ���)SYt[:fP;.W��Jh�|/�U;h&O�Ǣ*{�¯��௾��?����YM#���rd���V@���k�½r>?
�����Q���Z�+��Ju�&�G��+C�J_����|А;v��ԝ�)���+��=�Db���Xk�!�9|�>�'S~��5�F+��=�$P=a�-)�,����gI����C��榑�t+�5ܳ q���ԩn�F������	0L� �d�A�H ��?�� ��"������*�$�-8�S!��y�1���l��f���#�H)[���:��}�F�ܰ�e��L�9,����TM���=>�	�~����,���;�]V��9�$TJ2��1tvD=�8ԳsgW|��BI�$эb4���ځ-���}�&�CղD\�<��_cC��<x�_)V������`��j���m^�_�o�#o[�m�����ғ��O���a��w�91�8���De\�I�q��b��xp�l-ELb��$�%� PZ�ZZ���h�5��V�����F��8	`��ߜ�
�}�!�W��W f�F4��VB�	�u���}3b��Wl+�=�d�լ�b��נ�b�tx�:)��D�]��D����z����c˻C~�Z�=�𪚓��<�L8	��oW��<�w���hqi�V�U�$e*|�g<�\h!�0�{.� (���esy�|�Z�|[�8&��������