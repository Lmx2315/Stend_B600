XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��#���&��8省$���uk@{�/ZӘ�=�#�d._p_Iސ�jL�Ev4X���k<�L��w�MQp��/W�Ӎ�������THoV�t�)[f���J%|p���׹��x�$�f�h��\���?�>KUư3��Rٕ�j�'/e�SP�:�4��-4�ߚr<�N���yѴ����8L[&:^�E��ւN: �X�����a���H����n���/��Q�����&6E�RfPB�h�_���{����z/Ɩ�wT,���<e��b��&H���D=�+O5I�O������Cȩ�N���C�״SM�� ��,�H,�>l[����9�$��^�ځ�~��-��A�~B�7��=���7��g��b
Y{�v��F$�&����0����/�� \D͉�W��B(�NW����j?Y�b���,!��B!���*	������l�nƭ�D��6�XdY߅�~��_*��jj+v9�1H�k��RRv�GC�Jja�Ɋ m���"��.����UT_��6�.����!�C��>6_�ß��?�A�A;Lи)�� �n���|
��aO���o�[S����"y�_�c�Ts�� n��!1r�����dc5�G[[��Ng�*��ا�_�<D����v7sK�����ݢ�=6�Me�B-��`���Χoaa �j�8�����¯�p;�� z��X�9f�#�{�����BP�����V��w�΂ѱ�Ы�P��w;xF�c�#�kP�" �-XlxVHYEB    152e     580��*;>tV@&4�=�
5:�D..#ҝE��P|
>u�
τi��5W�ͣK�}�*'8?U�+����>î�j�zS���r�ɵM��O?���a��PVZ9��c��@�S�ߟ��9��=���y�b�y��i�Z�<��@:�Y�>9O[�b��jAQx�h�䣯��H*#'�`���8�/�}WGʻ�ٔ:�y:�}����~w��U��@(��E��|ޜ-y^7���Ew�C$m�'�d�:?L�V}��敥a?��=��M�6��u��XrY�~i%��_�0�^5���AGrh�Is�@�����1���s}v���\�a�L�Cw��w���5�]'C"�q���@$��@��E���H�
���By�ow�;��g�M4(8�./���E@PQ���q�/bk�;j���cv����G��h�JS���G�	�U�����"����R�t��3sm��NZl_�.tw[g��
'[~_<R�Ey�����wE&p�����UF��:���hoPE�2�ޡ������v�NlGS��v��U�RX��\h��{C��m��hgrK���Ǹ��͗�y��`q�߃��]�Mm�63��4�f؄�U�\!6���	�cB��|����i�9�a��l����wqt�n�y�]\MU��4�r-�K�{�96�M,4g���C�*Q�2ϜV������:�=4a��fl*B������>[��Wfq��A:��Ƴ������;������[I<k��c)I��e!�q3>�%U�����Q�N�o�Pʉo8ǴN�Z � �B[�'M�����,�����^m����Y_=�v�np4�^���L�i�N�X��ΛջH�� I��:s�.m:��m,u�b���m�{���7C����Z	���i��D�aD�z���JKa�dHKA��
 Χ�V�)GA�P:�X��Hɦ��#	e~�'��}{������+���c���tv�:��W\f��_�h�= ?�>b����*?�e�\,y1�K/T>�V�"�e1t+u.�����@݂U���N�y������/)��xRa�T���u1���V�"��
�[�X��#Y�~�?�2�)�ar����t�j�<�2��o`��P�~՚��ދ���zcae���N��6hm��]��$��9}5(��ĉ��ԙ#wYk��o�<���y�hVO�V£د�B����ty)��Q9�G��{��qn���)��D�8���(�͉	�+��{-;��r#B�}��Ҕi��E=`�Q2/��`��r�_"�XbV�&1�&��u��%5";�Z��<�"^g%s�@4i�J��: �vF��V�8���ø�?����?m
t�����'() G������_�w	���zpnm����j�