XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����w4n�I2
�,��K0A�=�	��	���2��v(�b.�G���d:���e�P�I���Xh��,ѫ�����n�SVKOJgJ�2#��:Ք�8߅�F}./�,�=�U�hٔ��������� �@�M����״�����t������cƛ33
�fT"�q��N�
��|��!PD<��]��A�.a�^��톁��u��������`���ōMX�Je�_�K_f�ɄG����B�S�n�40-i�3ۣ�O*��W�9��h	�L<������'�\�N(��oQ��á5j!�>�Qmj����h�C�#4���ʪ����r,����6��s\�k��2�� �dz=zz�Y�)α?������-M�IJ��]�gL�F��ѣ"��W�m��{��y3=y%���R�a���jD�\��ꠗe{��
��{"�~�V����0!� ����iy���a������cW��,���n�ζ�OjŖ����﹅��br����319-MF�'��O�������1�vh��P�z�dai���'u.I��~"��PȆ5N�p�������4�KV�b�"X�ƥ�3ft���E�Gk�6J~*G��z�V��H�V^~ظ:�3��K�R_%L�l��.���UB���Á�(����ǖ`��D�	ۮ��B�%�x(ӸO�X������a}���9��'Š%G�~~��j�y1�_�����=����E����f�w�]60V�4?��`��-���XlxVHYEB    3c92     900S�A�Z���2)|̖��*9�$�2֝�J�����On� '�:���,s���<�[}*��x��?z��Ʊ3Z�Y8�����X�,�)����>����B��Ao0Z�כkV(y�����^����ƅ�<�혋\aB�=�w�R~��=�$AvA��g8��@�� 	�n����A���䦶 HpKj Ô�3%�ۆiF�T�%^��+n�������^W��Q��R!n(��w&�L2�d�7��t�����XE���0b�r��]���7qSٵ}��Q��#s��xR��A9ٜ*�/Pz��(�DW���R�{��?Zp��P��ie�=�Q�d0�83��^S��ni�VPSu����,��̕#M���<�A�D^S�J�D��&������5���!�.o=!H�n���j�0�ҷK�re�	��..�apǰ�i�;#�MY�*�Z?�����}N���n���CO���VI��}�&�ge�ѐ�f�����?H��(m7KG����F����Q�l���xL�r�̝�_��R��5���EDk���5%y�n�v
��U��J��{���0�H�Hsl+� ��h�a�� �T;jiT.��n�<��Q	�vt\�p�*���<�n���V����
C��3r	��@�#7XY߰����BÍ�v�FD�Ao�1�ݟ�<c{�|�/!������Y8!�.���kk�4o��� �7-��c
�@ ��j�����:�sބwu|%���f�G�0a��`W����;AQ�C�><|��,��*I�b�&�΂"�3�E�f2M0?W�:�
ti^��krx1�m�nZ��0G��^~<
����֞-�C
��{�����?��x�v�ʊ�r���?�<���*��"!c�M��Ο���2�hAk�x���ȁ
����r��Qkd�czƠ's&6�C��ĸ�+���Gi��W���),R�n�S��5�y�y __�q	ѥ���@�����`p���}p˄3��KE����������FQ4��0���I-6I/���[|Hj�X(��ٚޏx=������e��]����������]~���u�_O����&gL�XJA���g&�����B��]q��{2��wWb��V��-�ɳ�!�d���h���}b|�і��y�c�+0����}�Z�lp|뷣5{ə������3Vڣ�Hs�D�-�=��M��!�]~f�4#��^N�JrAbwD֗��?
8ѻ�,ޝ�A?�Cs3sa�	��u8���*��hF�:`�S�W�9�S�J�� k�]u��x��}СS����e��	�/����Y�1����q�6�~�X�����i�p�����׸����};���%��c<����tx]���Lg�X�t3���P���4~�U�\�F#��eo�4U9]�4��=a�ӡ˧�<��1^N޻&�lg��4�V���8ٻ��%U��0�8�N�r�n�_9�C�G~�X�5+N��]���>c�����q�ן�ޥ�NAJ��B��ȵ��A�"��C��w���<��2�q����	j.\.����*�� ً�@�	Ѧ����v�Q�Q�ӳ�o�bi��⓶	5A�6)�63+&ŖXv~��I~`��)��3g?�ĥgX���J�d�)��-�z���{*��	��kN���a(y��ʃ�K����>�ؽI�!L���؃cu�d]V�a&��@A��	��:��]��搱�����q�5�U�r�j�;�u�T�-�qIpVa;�/�=\tG|�ũ����'�y�v�Jp�3�_{*�V�lf`;��m��l��p�íg���k+���)T���>Z�����%_B��\��Bqڬ2��d�'�rX�5�h�	��X]'����{�²lKP=.��A�2�BM�$�J�]��^K�J�Z,SR�kl���>�߼����S���w��BhÛ�g�c^?_�i�;�aH�!��8o�>��C�=�\�O��Kbͣ�;�x���1<�����llّ�w����c�9��&���w�/UL0<�'����{2ڲ����d�x0���ܲ"t(LO[ �3N���4���iN�����7�d���?� ��\�m_"����Sp;b`�v�����l���w�«L0�h͸�2+�����TA�f�9�F�L�Z~�o�����4z�5��i�/8�L�c[�H�X�pP��|�@8,�;�G�ݮv@n��H��B�gyp�l&�"�i��~�K'8��q��j�B(��w&G�ʑ