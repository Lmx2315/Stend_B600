XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���k�	ݏ.�jOu�d}�J;�Rqe��JI��_�����סh�\{t�/C�ۦ�]���:����# _��o�X�5�J�ǘ6i3h��e���۲�h�>��V)� �}��Y���+z��'2�����N�^2���Pm �HU#�n�)�	�]�"\��H'��	׀4����=���bP�9��ڱ�IA�/hZ�&����@�D�(X�d=��CjЯ[`�0)�g��U��h
[%���S~�H��V��`s��8��q�p>Ɍ��n>�%+A�h'~�?`J��m]��
�D1�|�>i} V�yNBU	K�K	�5����ǀ:��GK��@�l�g,5��E�s>�B9ƭS|�ǎ���?���%�i��(;�padw��h A-�kp�(e�c߁(�o��ˢ-����E�P�y C�/�'r�LT��5
����L��Q
]��o�m�'��8�8�7��G8m��?`�@� �����K ����(���s��E*F�'����x���뼫�r7�w���n?�H�~Z��E(Sц�E�t5�B�1�]������']���=Ұ�^N��ɹ[����A��{�#m�������CN];X�: �{K��y�q��$�nt`�����Oq�o�Md�r�l-pqq��x+&}�������p��/�i���>S���+��}B�@iR��m�Nݷ��Q��UhW{���Om	�L��{�É~��)`���v�w��\|Ӽ�	�>� �[K�`U�loXlxVHYEB    152d     580�.c�A��y�(N�ؑiv��$�Yw����,�0�i��dŧ����`/H�/�"�Г�M�xk	f}�̓�S/M�N�[�ƌB܇�㹞��Ϥ���i�ԯ=�\�楈��C.�G{{��CW���f�i����}<q��#�}�
���@W���*�D*�'u�n���Y�&/<`��::z��{����cC3�v����a�ɲ��gpZ���Ed�
U�\(&���F��}bB�|��W�YA��/��b�,�E�ɏ���`��i�-�7�E���Ȟ� ����'��LS�|�Dا��.1|h���@H��շV������D��dx|>3j�����h��o/1(��U$5g��Uk��E�'LDB�L��HI�9�Ot�m�wa��#�����D�D�_���}t�y��M�e|��s[���kia8�O�=���'���.y:�s���Lj���b����	���Wi py���Õ���L����*������!U��6;!����-��)y]�[1:��ϡ���܅�I|$3v��Y|An�w����1hG�9S��q6�\����z`�U�<�F�����_H��m���hJ��<\Qv�ӫ``��E��@�<o�lO��s�s��qWov�Ukd���O�5�P��R�t$�#��V;4�V�:��f�ފ�DU�;���@�f�3���=�k��URէ0~�I������F~>Ž�h����ΞAt^ĺ��3i-�{Z�qxVA�'�Qvs�g����X�,1����֭4v2L�Wٖ=�gzzpVh�Ef��pP�/^)��j=y���M�-f��{>�yi-?仌���K������4�YX�]�ޤ�,��I��n�aK�#yQ���C�eዱ�������N)T��D��p�����w���խ��Z�9�7���a����~e�8���7׭fS��9[�lu��5͜���`�����|�|φ����3a�q�}��=p��,��I|�u�mkשr�ućI4���L�s,!��,�wo���X5���?��D�V:Xi�)�~�����z�(�@��vPG�uk�.<K ���M����q��R�ɘ���qʭ�/;!s�WM��GF�^jܓf�1�5H�'C�_���>���)�W���g����yL��T*�|�ť7=����Byg�D����x���a�>I���P}��H��]#���a�yG�[���ts̻-E�_ಯ �u}�E�XcH~5�n�D?$�|���J�
W @����vpx�r� �Bɻ{c0��:7g�Ȝų6ˇh� Gb'�7��^�����B���`;B4J*o.�xKJ�rT�8����q�?.4���wj�y�4��T���Ie-�t~�xK����%�Ս��ߩ�