XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������{���\�����/�otO��K��︴R�y��.��:��8l��xwP=��G��K�t>��8�x�ї��(+h#�[0O��B
�C�G�z�����x�7O(���v� ��y�XA?�䦼iͪ3�X��;�Ue[D�W���ŷ���Y�*�n��f���ș.S*��w8�����Ba�*-n]�Y>�q�ӆھW��	Q�6�ڋ&��R��(q�xny@G�D2b�:����z�D$WvԤX�|�SY�Q��
4��ĺP,�i�.�񖕢�@.��d����{
���������-Jk~+l���]�o�/�t���<!����Z42���S���=��O��h�*u�s����Ԁ��Zx�<����3�m�"v��R_0�T��|/�%�ea�1�F�ȃ�.�FD��]��2ǎ/���2�F�s��8��5GoY��?w$������4���6��8ds�ujnV8�Ps�Y~���eF�����<VWX��bOX���w͒���܈�{���it�~�*��&HaO��^e"�6i�R̂�zE��V��ޭ�������q^Q����"{fm6��7�֦%mW�Ca��1�B3cZ�n��O,с���Z���iI\�-=mz�t���yv�����O�7O��� ����Ҁ�7�=��u���[I8	feap��=��|��h�� ��p��}�wR��>�xgO�$_�v���T�7!��8]�C
3���S(�aQ6�K���@8E)�XlxVHYEB    3c8e     900>G� qK��o4:/�PӘR�ҔX[F��o/LF`XJq��3�'�x9�����~�@�&�ZU����z�̃~E?�h���L��#t��}��f���8k�?��P��`k�E�F�����%��ȉ�R�cݬ�عu�aY��B�����4��l�C�QRM�S?�'�Â�vhB��+3��!W�0�_Y=F'�"H�����S�V�F�W���s����]9��a����_��Dn��$���g�+y:&�x������zS#�_�0��$k��Ap5
��O6�#�CZ@����Y�W�q�g�Ly�Ь 6�}��%�jVh_l��D]8�yBj�F�'�U���oz���78݄Z��?mf����q��<�v3S��6��	ʾ$[d0+Z���y�@�c��2T�"�����'�-,_8�h�[B:�d<��-Pwu�E�(���`D��j���ɠ�Ɓ�I�eTU�2p8v29�S��%�8���!�3;(F���Y��f�ء�}j.��X�6K\j��͂g����F��dv1amx�!���b�74���-��|Fc�aQ0W*�|��t�4�*��\���2�=Gw��A��Ȣ�v��vwy����c�^���H�z�C�#I�	֠!g�}�g{;kA��7V�n�)�h���W�L�iH�4��P�%H��>��z�+�D��f��˿�λ|ȠT0�լ��Lx�55, >�������y(P��fI���f�U~<��[?�X��'�P���BE����'̐*�3I�UQ���Q���A�l,{���c��ʈ��@���ڻ@��/��3j��N�������c� ���i�wFhc�Y�jR�]Q�y9��l��vA-�"�[�۫��<�Q��yC��0��Hs,}A��)�/n�6{4�vԵ �Q��R�Bx���@���e- ."��������e�� ����X�q��y�ε!�WrXm�=9��"�.�-�Y.��f*������jt���ab,��H�3;�E@&��Ti���i��	���W6?p�[�E��;>�� c�1�KG��%0�@�X]��S/��e�Gކ�[�qp�G�v`��`��}�?��O��ue�l	z����]�{�4$Ts͸��1�^�K�X�Ż	��K�t��h~$G*�o�
�`�t�X�I�K�\���R�/B�2�{x��6�d�!ij�sJn[�(���{��} �b���ք��y0��+c]T��`n����뜣����bLDOd4�̹&�s���	*��ߙ-�p�|[G��'g[]I�w��\�;�P��9TqH�;=�L���������į�BcM��`�X�V��вK�M��ztPb��|�H���$�&��RVY�Ģ�����N�v%��Q�n�'c��s#=�<��	��2/!��[=$�c�#c��/�ZQ<��ӥ�bp]���2�..�g�2��<s�ȅxH�x0[T`�4�2ߌ�B|�m�����ds������E�����/|(�#9<*�N1p�џ�OQ�)/��g�,v�Y7�X�p�5K|��s6�P����e[,��7$�� �]H.0�c4�\����n�F��5�u1���b�/�pN����.l�ܽ��(��]�=Oc���HN8ؠ��o�I����5�^�|�U�v5D��1Fv{�'WJ�;�}�[�"7N��ѓj?at��h���H^�.UW3��E��*�[�jdV6��R�vJ��6��ǂ\6(�4�6�4�2��yb	��;�}��&�Y	�4	����ؼBx�l�&����*k��
�\˦����֩
t#����؄�e���?&S3�q��� vii��|����j7t��TBR�1v����ԡW#@�'K3BC��z�:aR!�s�7�F�%�0�����,�F���Wԋٝ�2�[v�/�Rsk����'�އ���[?Xe�:��\
�q���(�uc�*;a�' ӃP)#o4,� �����A�%�͟N��;�ȑ��B꒳w/�c��W+� xLNC�"k��N���^<t��"�\v7��v)�>���s��C��7����U.�q��� �[��x�U�R�<m3�WV�9�Q��2/9���YOm5{>�a�s�� ��ĝ�D��� 	��VbL�|y#u6L�W77�_00�`	��w�f�q1�I�ZbM9��GlZ?@�s�7 3þ�52�=�ǟ
(�D�7�]$�jp���<��l�&��>���+��QT>F�W��T]�L����#k��|��~un����<�