XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����$':J��8&���I�8`.�w窇��ಬ�k�Ң�g_����w���5³���d�f/��%�Cل2n�zX����#���%�}���$I�6(�F#9��HNj�404y;��{F�᭔���=�H9�^��Ҫ,�G��~.4"n����`b��wgCês���j��h�j��(����x_�	�Y�6���	�b��p	�2��}"+%hK��O��y��e't�`��h33���J�
�{I5۵�'2�&�݀$P9�mw�YT����r���v�Ȋ�Y�$|��=N-Q	dXQ�C	�>Ҧa&!	G�x�[p��f _�*�R���^�H�9�lR�4�b�4j�-����XM�>�n�7�w.���-�]�8�;5V�'b8e˂�wY!1&������h��`�n�gMARU�/��>k�YbL;�u�.��:%O���
5L��]kbeo�L�ws����n?]ٸW+:+�`�Q����4�SY���.���F��e�R�d�B��u���p��/>S��<d�X*�� v���' ]O���bb�%Z���`�<�
���WpT-���qC�ё0]wLD�߽��>�X������F |1%�{�ϝ�4Q��9@رy�8k @:�:�*]RJ�x���d=�<����z��2�a`��4�/�5��kpN
�ad^��/}l��e�_ ��/o��v��b/$~���3u`��>�^ �f ϖ��`�)S�
7����Q~/�5Ѝ��XlxVHYEB    6fd8     c30��c8��QJL]���k����r�y�y��X�گd�hfhM�]�H�+�B�:��� ��]����')W`#�3Xx�2g�65
��"�2�Y���b\)`���c��G�_��a��ؐ�>*��C���f�7��R�;X*h�u�*�	����z�Ao�0mk�67��C�E��'z���޺��{[۫��ݐ��|x�rJ��ܣn���K�t��;%-����>]I��P�*Za%�$��y�n}l�-���VfZN��%�*��AtC�0Ɣ��֟Ʉ0#�N�N���7���%nS��H��I�^?�Tq���7���� �:L��ƞ�N�>��
�y��y�SQtl�U�fJ���a�^�]�/��U��ydU� d��zASؒ�z���AF��rA����Y)�6u�%����XW����\�E}���{��R��q�� nM�����)����(�{���^�8f��+9ȗޕ�'6w�J������-h�^�t��޸��C�3��\:��w�p꤮�L�Z~�ݝ6\C��pS���͹���~�q�S/y�W����Э\R%�z*��u���C/r�h��t��g�)d�����1|�.�=�{�~p?��`ǉJYh�Rd���dO1iMg��3�]`��=�]W���| ��&�����}���̖�v���U��Y�[�M�T�[��q۫���`��[J��Sy6�T=��/��x�_�^ ��sz �ڮ��������IpW�����4�B�=g��{�X}N�d�H�$X�n�iA�ڰ�bg�a�bCz�̥�FT�^�qS��|��/�p�����G1�a�8���\�\���wN�Ѡ*D{B�X�"Z�If(�� ;�����@5s%/�+�)��[���ȁf�����"m�/�gvГ�����Ae�`D��j��c��8��]�hzS���4Bѥ-��cZ(�/���Y$��k�����ŸMd�dʩ�H��%�/Q��d�m	���Ҿ�r��*|� �A,*笺���!@��ԈX"y�"��[�G�ma��T��[m������Os����c�0�#?��	;��L4^0��fR2��V4�����%=؃a�,� #��Ћ�+E}�N��
z�3�l�O(�vs�����* ?�QM�@}9?���yn[�Q�*�ފlَ5^�c��X��vce�����q��M>H1�^	�S����`
�@�a���@�� �����6����9�5G[�*ɵ�tT�ۆ��1��JՐ�d{�#��>G���5�N���oD_.�YS�]']�VE�Y��S�-�/f }��y�����?���D����L��Z���� ���Ib��6��O�W�b�u,������h�}�䈰r�?o��$�?
a"�֋8I���������G�h��s��I�6����#��l���Ĝ?{�koF��8����`�%d�6XI�����2��,3���=��;�8B�+P&4�;$�.���b��S�ȅ�XG��1����Z>��N6����%7���*p�~ @��,��5�b��^���l�	��F �%U��U#��B��P��0�?�;�!^]���<�<R�FW�'� �[��2
;f�ghD��_�p���I/P��a�d\�������Mxbu���I 8V~�^��1�)p^��dX4~qܣH��wH��E �@����g-��K�T
+"�Q�1yQ�uL�y�/}h�r���9��'a��v�e��2!T������8c6t�� x�\��� 9��>
u;�Q��O9ߍ l"e*���\pz�K�D�G�eY$L�(YL6��^P>A$_|,��a�"2�6L\���ni�\�#B?a�8)����I�E;���~5�p�m����7�*��~�l #ւJ,aA ́dժ�-��q��O.@��ip��҆�N�xѓ��J�ʦ�#mU_�p�l�
�H+x��@����m�\����	<��8�7$�p*�II�E�Z&�3���7��:��ޑfM�4��K���H�8b�UkGE��68��W� �*�O����]��4�$C��x� v2T�e�P5�=�����d�"��3}^��)hu�͔�Ԭ������}�SZ�f,{����.��2Wy�}X�-�}L��p!����0�_K��Щ����Meua������*|%K35ÊM�e����z;�m��/��{��4tR��_�3q�*c\�˖��G�
5��n;g+�*�[ɿu�������w�QL�!���h��,6���W-�-G��&a�?tg���ՁH�o� �@�(Ђ
.����x5��`H�JC\>�.�}�O��n��ԏ_�h�<*N�	������$�'��,�YgJ&d�>ߠ��VT�4���ɶV���N�(H��ϵ�L+V�\�������Q!�=�[����G�l��'�C�jP�]��s<\��KYH�t	
����x����	X���.�rh�[�M9���X�T�M!2�fY���� �Z`��S��; .!4-���jgR�A�_!��C-���o�C���B�m����~Fw�4��J��38�uN��-XGzv��b�� � ?6\��`M��F���5�I@��.���0:��Y�X�I[9$R�n�}�낋Q@Հ]9�c�"Ǳ� )R�g��j,���iN �t�0^W ����(N}�Bl�@�G|z;d��E��o+xedӤ�)O#ZS�RO��jf㈵_(�N�����U��`��h�=!+r8H�S�LgP��ִſ�'YZ�`�
PC��nh$B���z�&�9Ԓ�#�aV{p�\7G���S����!��o!�&�i�f�����?���}%G7�eۑ����>�x�^�Y��.8�3v0D�?'/ m�}7k�5��#T^'2�z�*h�J��m`�Hޔ��HX����J�u�|	�Ͼ:itZ3#�OhT!C+'�y���+�Ճ���tM��BkJ��
A�0?M�9%�;3x�9�k��f�ƗB��$wm����m����F����荆 (de��F�Z���\	�����&�i�k�0̈�z�G�