XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��N�8BY�Lܲ%e��~�o�a(�hL�ͯP�Oa��Tp�e'd<PXA �"�h�.'%�zx#i� ѵh_7�������r�0��+��E���jƔ\���2v�Q]���`�a5Qtʮy�fQs����`��P>�ևh�Eh��)0�����4s�z�F�sab�#�qpP^ͩ�_�?��|&y�΂mƋ(���-w�L��/VIee������]��:o�Py��u�VoS��v>��{��Y�_|����`��U���:5?��܅�8ڙ�ܵ�mav$��uO�evs
��d
%:$A��P�Of�N�!���|����՟,�Db�ǆ���� �D��xL�c�������]S,�ԍ��P�"�|Z��7���66��� �:�󞰷@�n��1�����Oz�s�J:2Δ�����D3�Pkt��8�k�"�̫t�,X���]�{/������K�n���Z4��#rY	��ț�(gG��������+���� ��rK4��B0�|�2�)�ȉ��@�6~P�ȳZ۠��X/�H�<���:Wٲc�Dl�"�r�n��U�?G�Pg�V3ey�ǜ) 	�6����y��I�hiG�����5�32x#y�Z��g<�k7;`泔,�齷����!���z#�&bx:��U�S���>e�8��<I��qΝ�?�����N�"I?·�*����=]���CPe�^|��ϖ��!��	�*��&���ye��u�4�������V��1��XlxVHYEB    fa00    1960���7���Q���Ю٭$�}�J
q��q2���EN��5֌sH��<^2����v��xw4����U�sh2��8Fy�9\��_t���<�5��\�^R�,k�^f� ��p) ���%#
b�ރ���~���~M�&XJ�9(�.�H��t3�k&�33So
�l�>��)�5k��-�N�>�4�ꠓ��^vl�B��xxoO B5qU�!n�y.��L��QU�$��(r�ˠ��~��I�Zl����Ӣ�� 4�{"I�.o,��t�z��vu��l�v�fR1^X���{z��M�Im$J b��6a) 	&a%YJɺ�<q�zU��)K���H����p�^��r���O���U�S�صq�ܮ����[,8�p85,[��s�1�P~��[���lwP��#A6\U��t;��W�}k'����#�Kt��� �:�N��ҙQ�闑M'�=���皣>5��+"0<Xb�4n��D]�aO��A�Ԝ�b'�Տ�}���\�4 �~LP� ;��0��ڡ���nh}\-��{����.�n��}��z�<���8�Ӑ+7�] �@V�g��B�W
�#~�k-:!I��z��jq`��E����?�/��z����2�ɔ�V��#v#���Z��x0�Ҏ-�_&� �b��4kf���.���w�������N�+��Jf�m[%KLF2T�$7A�� �R�L�ǫS��(|Qa�qkы�.0������%�S�[� �UF97�_(��JAt�7�3ل�N	HXqW3�,٠�#}WT��ug�����GU��o��p;�́:��_�f�9翅��}2<�"�Aٓ�ʖ�²��@u�Q�TZ�nW��{��"�4S+~�}h��5�%�#�[[�T+�%�L�D�k�OS~XB�w��~.����q��=	Д�0ن������3�4M+�J�M�.��rXXP~�!QL�ɟ},s���k�ʨ��r�{��� ����x�84[0
���e�h���$�)�� �?�_��,][��C���h_( ��l	mx�ݐq�Idp/5���2x�(���">���ސ�����}pc!c��`��
���j�t[ӖY6���s[���k |��g�Hff90�d/�eX
^���Xt<�|��gۄ/��͌����y�%YI�9�p����ۂo��r�������M�J��)�a��H�&���6�)����Jnk�������.U:Vr�Q�,Y?D<�K�m�|�m�JhK�D��X� %l 9���rܰ6�����UJ����/S�}����s�~B۠����U,=du޻��:��\���"��Z;Zc�}j��{5�D@ΊeƲ(�+�ӏ.��^?x��%�kތ�Y��i?��)�[\�����������?�n���>��c�Ag���5�u�a�1b��Φmm����ڿ���$,E%��u���J:X|��������DR�`���#ip<X��� �p�;��.�����ʖ���*KJ*(:E�|�K?7Y��T�׮ɦ`��2e:��7��-�;JS���q��Q���+=��y���lg>}�7%�Qg����Q>X�^�K9�cws9V%,c}�@����MF����c\�)�эW��)!�(������i��	4GMo�CP QP�*.�Q�;��+9�<����$���R.����YZ��R�f�3\�&�m{7�"3
�;�����;�ԅ�e���]�����Og@�V�F8�sv���5Dv�H�\�P���o}-��-A�P
q����|��T8�v�tb�rCtP����JK��=W=z�ы})]��`6_aL�X�U�8�}�y��|OB�^kwM�I?�%NWϨ�-�|��mr��)�W9�N}l'��u�>� �'ҁ?n�xc�9�I|�ގa��RR���˻��z��8���X���:Z>dP����}�ka\�o�}v���j�z�a��|���4 զ>�*e
���ٙ#�I�4�5��R #<��G�(��,����鿳񺦠���9Zl��I~�2���
�GFg�!`T!!�AR��6��A�W��ԟ��]weO��qz��`jW6F;B�\+����3iŶ�GNx=��Ip]�b/r6��B8+�>��V?���,R��l��j��AU�O�Ap_<��k�D�%���6�K3�My�f.�2���D.�Z=ür�1��7a�D����
:A�e��1~s֙h���>����н��(a�E0�#S�#�cu��8���x
hD���\�͋�F��W�.�'��s`{,�5�L�p�Q"�@�������2΋�N�<�W��[jZ��%�;T�1?�S�y=T���y^�����J�UA����l��z.�ǈ��鉤/��WeZ9��;�,�a����[�(�!/u�ުEL˨��Y�{�<���LAQ!֪괇 ��Z>iG�/��͹^�u�	���2��p�S�J�EȀ��m�8-?'����8$"�$V�njQ�P+��5`�e����6 4�u"n�ō����.���$�y� =��Lw����!x[���~�nkZ�yC���/����~\r��h��TE8��f�f���(�s8��6��3qѢ&y�H?���l�2˺�!�g�`�+c�����T���O˪�1���-��)�[�YtB�e:KX��Y���9�$;#�vv�K�	�l
���������pM�����Z�N)[�?z{�[xO�J��F^B��
v�؝L�n�����!�ླ�ʝ�_�0�@|\Dү��/�*�Ju�/�=9�,�lfcH�{�h�	��r��&5���	���`�*����T�ɠ&��&�Rwp����fI�x9 B��!L�9�TR����$wPP~n�D�#<�� ���Q��;�{�(���F�����{(le7��������I�L)'�� r1,p�(x����%0O>�%�.�U��[�m�4�g$N��Dr�棧{O�|�<��a�⸳r���GTt�Q�x
��̙d�G@L�K������ZU��!66 ��(����N�<��Z�D�d�%I��b*"/�E�/� ����݇�i��S���|�t�e����a�3��ͭ }���BN�I���Z!DLߛ ��s��1\)7�T���a6�wd͊i���2�Bz��풆� �28e��*�$�;Pjȳ͂`=�%`���t!c�?�bze��
P�Iēr�߬����i��/��{�Œ�
}��(�k<�W&w�&zJ��&:��oL�n��%����*��O(b���~x܇��楟��9hNҩCZ�3������&��c�j�[z����͙N �0�ג��tr{D)de�m%�B��;��lF��P.n���\��Lx��!���r�|���P)6.N�U3OWX��BE��3���@�(C�eNB᭩|_�R��ה��w/^tl��c�fs�5��G�s0���{<���Wsc/�p50~B�'�0�B�)�8�˳x�]}F(�Xw�h����ت���q�+��11��[�<H����c�6���n��]��S�L^��9�])a U+K�o�Cv���U�LW �>]{z�}n&�c�%k{=����RfD1���e��K��L�<[��k K�� ��p�d�g'����}\|���s��D՜��(&A��#�񁔡��[��I
�CO�Ey��3ICH#@�����މ  �L�	0;p�)m��V&$�8*s<;9L� ��|�JY �RZ��q�y�P1��sjA�9��R�-�KBa���Cչ�����7�Q\��?C�_pC���w	�@��JN�R�W#�x�[�<��Q�sb���������8���ޮ��.�9H6�7����x
$)f<�J�x淀9�J��>��[%����0r����1P��cKP�W�7�rD�\?�����*U�39Qmy�8�N@�%f�7��9��8�{>�=mD4�T?�S���
�ِ�5be���P�Kh����!���ⅾQ: d��@D2BE)���@m���
�1ė؉_�4P�ҜF�=	�U��3A�=��P�U-�D�]\@*�Z����A��J�����ĸ<�&D�o�,�S����O�9�X�>�S����2��z1�}ւݐԑ��ʹb�\y�Oz�/��>�a�h�8�89|^��ل^o.Tm��S��|X�V��LH/U����!i�$d��JU=�/�(�p��n��!��X� D�׌�*��V�Ѯ�;`(t�}Rh���E捱m�<�D�ͻ���EDݤ?���g6H�B���c�)�u�ˇ��5<���l)�$���"TX5�=��_6�^1��l���[��2�*J4,]���Q�tݭ#ۻc[��h�:�ZW|+���?��S�0��0���#��/Ǚ4ژ
�Ik4"(m�.��b�B\&cD��Y�3���aR�dc Z��4��8EV��"`�@R6�ͧ6	�B�N�KO��?����+F��DT?�Z��t(a�ٴ�hg�Ik, �>���2-T�#����K/fn��\9Az+�bw�'��Em6H?9��Z�X��<5l���?=y��4��3����U���a�/%�ttg�x�8��w��}$/u�4� �y?E7gs�!�K��AW���SN���(N6F����J�w]�5�ՒvD����FTY*�V:���Н<d�F��E]�-ozz d�����K����ZZe�QnPN��MCW�n�7�"�8�))�����Wث{3�Q��-`�k]�@�{����62��4�OE�X���~P�9$ߍ���o�o'��\�(���>	��������$G5;��e��N��KQ������#�7��n��7݀�j���6�mS��,3
�/�����92�Wh)��H,�L��<2[·�����7��z�q���0l��0L�׎بNx�+�m�-��5�XC�X<}���OBGs\��~�(��°*��p����D��*g.J��ѮF˔�Y��h$+9\{ԟ�(Z��0�:�f��4�*�|���NgɫG��-�A��ƌ���2�B�J=:d�G�����4܌H��zRU�|-��^�
�ό�|��P�u�O�.~��\ń���kަb�=�����m;��D�
h���%������2^�m��Ǌ�{C���{�~��2�Ď$��D��[p�"�̥IM�L�Q�mM�0.��������lT��I�+�K���O�$�����_����[D��' ���B��������~�Գ�09��?��:8�O�m�|�{�a3���Y1�B��~�% u�"o?��V f2��}��uN�z�S�+�0��4 �m�"R�X�*�&1�Վw]"=�mIJ�����W���Y�ܝ;��m�����*����:�v�<����+h��9zHw�*���뉷<���d4[�����@�Uu׬Y�B����ֳ�N����=h� ��K���ٛ��_�[�X�p?��H9�<Tŗq�^��q������~hM��0c��	�"���U�0j\}c�I͂�Dh>�agK�rJ:.�.Q��خ�3�D>�	S��l_�i�^4r�!U�t|����fu�S1��Rx��Q�����߾�kX8�ټɱﻚ� I�f����ɕVc��A���E�nٚv���-��#��ॸ�B��_��+�vw��E�r_h�3�L��^/�E�[R��#�&��x$��8��w�{�
֑���to��$�F���qy��ox)D�?��x���2���	���u���9D#N�O��'��]�I�j	�++�_���9 ��m@�3����/2������n�+�;9.���2׹h�/}�՟������Jm��es����z��j!���ѕ��Ȥ��ʓ��ֵ�f�P�-��|��u��q�fRn��pwN��V���o$u��j��qt ��~R'ǖ��&���qa�M�x�wP(��w,�r����|�?�?��h�'��TӳXP��PU�����W����7�}D�@=>M�wk���Ӓ���T:q/-����/��m_��	�����,=��3M�������T!�m�K^e_���QO��?���!J��w��ѭ%�B�}�E�¶>��O�7r�]��M�t��1]��;����Cc.ua2�K��
���7�1Zy��NR5�Y�=��%&O����'�A��WL&�n�'oĦB��~;�e�pz���]�����ӷ}I�6��r}���������F֮�� M��)�����Vy F$+菿�G��Lܔ�@��@\(��3�dB����J�z�o�,�c��,�{�V��F������\���G׍�q����V�[�mXlxVHYEB    fa00    15b0?7��|Y;��`N��9��-���:C�� �W��^f���H��F��	�9h2b(0?��u���cЦ����^�i��bd)��Ջ�r�MF[�]�&Jm|h@�[�O���X�*ôv���t'^����)xlL��jGk6]��he��58�b��ה�~��]ĨN�߇:��h.,���m�$v��a8�:�(tw�W��"^e�����`�_#���yOd4^�mg^����d�W�l��oxV�EUE{�\�Ֆ-ݳ[x�Ns'�g�Z��dx��]��A��yr��Xj��D�84P�׾N��.��1�|b1z�� ��m�UeŶlA��"���B�[�!#A�(W����<����hC����,1��m;@���ӭm4���pa&"���z:΄`��	{�D��ם(l������O1T������=S5N�U�X4���%�1�q� ��Ɍf�Ը�,�2c��~I��Vi(dC�Z�q:(��w�5=���O0�c���ސ�fY�s����l��?���Q�6��"E�Ȫb�Y\e���7�I22n;�L~H�I0�T����I/Ŧk]�����(F��(��F�V�,���cQ���|�ͪ�0~N�g!��+��l�����
֭߻�m������&>{��L�A�e� �F1v_��-�_ü/�B�0%<����[X����	ޙঐ�oz������>*��ۥ#}C<��m�y]/7j;F0��=̠aڒ| U_�1	���%�%�]�(ĵ��
Ŵ?3�$tg�\�&x9�O��j_�9u�O
p�C��[�/�
'�W.>���캦�ر � �wn��XI%R�F*LC饤�d�ͮ���͹5�p:��H�Z{_�{d��f�$�($8�a��H2�J���ڿ!H�C�k�'9x�;�%���l�G"��'M�82��ϊ�G�Cx_���[��hӲ_	[������5c��6��ߺ�8�chƇƩ��b6��
��F����z����T�8�%Tk1�"S��%�h�.�|�<�L�Ò��m�!�i��9��%�7&�����i��%ǩzm�Q�Ǿ��������'���D|!8D��X�\L Oz�=MO�cn��u�fٚ\uA�o.Ɣ���=V��9��l��]�B�W▱�/K���-��Zg&s���݌t�ӌ6L��+�� u2d��V�YqvTt�	3�ȁ�i��$.��b�?�i�5����Ű�\��\O.�}Wݓ98���fe�O�l���0r���	ܳPe��Z[�#�l�ksTpp�9�A��'�vG�cE�S$��Y'��o?��^����}�y�a�O�A6�� �kT�ë�cث�
BЅ��*�XZs[*��`7y�^g��R����;��O�W�NY�<����<�I¸H�o��uBϿ���:��~�Y�͹^B���c0$���!�]������9������]���$eO�I˰�ym��c'0�׻A@�S�jD(� ���̫�x�*@krTFS	".r��D�D�ɿfi�^g��G0ꌻ|�ތ5+7A��U�]KG3�(ـY�N��}}K�Zu����qXK�6���w����L����u�h���q��h��!.�UR�gIk�6x��c2�Ne��]}�u���*_�s�ѩ�0Ipq����\�� #{��ƈ� ���WVq2�3��Ȁ~QgdOCj&h���Ԭ�o���xyUS��݊M1Gz�q��y4�Ⱦ��ݝ0��<y�$,����"��%�m�)x0\����]�����]��%.��0��B�Ϡ¿���������^��c��
���>�@�/l��W0�:��6���j?�{]EJ�Ư$d�d-7�L4<�s0R5|�E���^���+E>�{�r�q��&���?�x<bs��P2���cN?V`��&�!��Ӏ)����YT�!�֚˅w�j�X"��%��J"��&�v6���@����Pou/'Y'Q�K_�MP�D��h���u#W��_|y��^}��`_�����n��W/���pR���4�|o�Ө2�n5�uGg1�`_�pT�����̏p���S|!(����;�J���C�I@������6���@	�{�1hF*S��Я��V+�:��QsFV%HNy�trc4==uC���>:Mɐe������͢�z
W/�Kp�Y1!
����Q&��n��$�x\��ʣ����g��į_b2M�N]-*������˔�SQA�py �+C!f�̧�F�"�ܣY{X�]�ۻ�(tq �#/ۡ!��(�%̤3����A�O!����w�O[ƙ�z�#��r%��� ,��Ff0�'��%dD�Qt'6S�g�(>�気��4�rK�; ��HQ����f�jm�g�� 8N��<$Z�nٌ�go������Z"�K(,��H�]9�y��>���p&�l5�a�}¥i���m�ŧ��?���s�����]q(#��޽�	n����7a{!=�V�z/�)��P�=�"	�1\��B��g�,����"���a]"��߲n�s؏���6ό(����S�1t	X��0P�(�
��t-.�(r��<�R,=�@2�2��V�B�<�E8ɀ���ku�a��f�-��~�R?�gm�zt2�*������&��#����]�p���qu �F�e�����)�G�I��7{;�Pσ���,�Sn[#D��!7�U�L˦j�&޼���Ў�s05'>��?���?g,��� �&��83�I��;��͎��3�t�?�/{�+�ᚱ"J��屉���3��i�$�M���(߯�8|��aq��I@[���gO��G�6~@�����-ԥ�� m����9��fc��A�Hi1,w�1�x�`t2��X��4;.x�]+2�<hl�H�Xd5a�ڵ�DhzR�h`�hy6{
k���X�db��K 1~�G����g;3c'm�c&���S<�������7�Mt���M8����2�� �I x�j��7�I�UrΊ��� 9&�p�qY!8���z@��},*˔�d"z�7��G1ϛ���vq���.~��;��w�i3�´�=���wg1�J1NB؛ZuJv3.ܽ7�'����r��"��5c��Q��x|<g^Z����yi�"��{�P�������J[ƶ)���Y�r
d[�̓�Y�`�ܵĖni���J�1��*&|3�Ef�A�����$�zad��BӠ<�x��g�8j��&���ȁ-��T���)8�E��Ft�׶��f����jː��F
[>ծ��Աug�{��g L�I(��V�$�J�4�*�
i:?����b �O6%s#�������8��M1	&�铇�wu�������O�q=lI�2��Q���*�I��b|5�x�W�|^�,�]���`!m��^���`D{�3��!ao�;�Ə��k�#�P)�\-�:���h�q��������Y�h��+����x}5�Qy�6j�	�f���v���(y ��	{�}F<��1m%�,b&D�l6-����ߋkϏS�NA��4lYVXHaVY�|���t�^0�!��_x"�Y�b���ę�s�^&�/1���)��#+B*��a�J,�~a�[ź�s�Xv�A�ɉV����.JӞã���X�-f��_
���g���M�ĒYX�)���Giu��ڸPIn�����at�	ߕ�0�mD������BX2��:J�[�)��G�1�2{ik��� ��̷ٺ�k�*#l�hI��d�}ً�a ����;X��.��3�J��WK��:��=]�I�D:��P��&~��x5s~�������o�t~��"��6x��'5�ߦo��A]�ƈ�G�����1�c 
�$��?��wo-�ׅĀ%�Jg��>�9.]�md4��Q=�ӷ/��t�c��;��l���_���0y��3��@k3�G���aV��L�p��
�@dAN�CW��Yxf���W]�i
�0~�vڛ�Z���� a^fo�<�J��I�"	�ҬN�V�b�Tc� ���^`&��·'y�ZX�0�RP��b��@��b$d�O,�F¸�Uy��VY�<��00m6P���%�)^-9������o,a�D�%XwJP<�9���ތ��~S;�o�ҁ-�EQ3�_:���_��}>�<��G�t��3	'yjEwy��O�A^NdS	<��-�Tq��������0�~NX�'N�U���b�☌�e��6�ܚ{���ňQe�d�sDb��nƓS���b��p��nGj��?%�a�f
v���?�D���A�ͮ��3b��S�r�_��z��n�dK���L��>�ʍc�U�"�tlkMw|���V	)�/��z��"_"����=�������e/d����5�-�5�|r��[�:b*3�����g��8-V� o\���g<�R��"!�����������=M͖?:Uѝ2n�Q#H�=7��{�� ����	��2��;�y{���F�z#Ǉ����'��h@2q�cU����F��幻P���R�й�g0j�A		��u��v6A����CۣJ��jc)*�Fn��X�����*u�����rMu����N��r�MQ*2ȝ) ���������E��~T��A�.;�!�h�d	�Ů��d]a_���I�nQ,B«?�${���YK������fR�b���Q��bi��5�3�_!^�yև�sV!p!x��k� OUC �3Sa�o/���~--�VD�5Ԟ�L��YC��R�*�ڲB����O�>��y/����*�5P�;����d d����߽;��3�oa��bR�~�+O�a���8�~��tNvpS�߯�q� BјYGU��q�ͮ)^�M�R[��X��)�ᘲ��:ޒ5�@a�:�%{�t��O������,�	r�(!���޿��Zv�
KJP3C���v���qtK!�.���L����ǻ�@�L¶���dP��\ޮ!n���I>V��������?�G�S�k2V�ދK\W��n�`u��σ_�I��G�J���-�Vd�I+*���$J(�����h���L���Tz���"�)y͒]9��g(DO#rv��C"@�����$7IH�k3@x���zS���<��Z�vY�ܾ�G�!V|O>�O?��`N��2��K	D�+j8����1ܜ1���0���<�z.����p����
K��~I^���� ��nL�푢�X�^ݗ�/et����t��42�/�Q��m(�p&�Rٺ��K���U�D���fX ���>W<~��顮����r@Lt��l[�w������4�"�������a]EKr�z~�T/f \�įS5ݸ�lD�N;�j�����=x�4��>�x7�O^�Q��}Y�9��3 k����$W	��K�t�`.0���m�R�1���k�˃ ��MJ
�;���޳]b'jXlxVHYEB    fa00    1600+�>�7V��[�&Vw"�7����8�������e�ڿ���XJ�`�����&G%!:�:z���L&�V��Q0�U�I�)�&'����,�G���ab,����p�;�����_e]�*�E6��m�#o[#e lf�֪����ED	ȁR�0!�8�1�W|��P߰�t�B�B%{��\3c�J�ۘC��A\_I���>��0=Sq��\�l3#�c �D�n��ޘ�����������Ҟ��K�g��ê�� �y�����M�\�ax4�ڝ7��N�,�C��Z�m�Ĉ+sڭ��iC)E�C	`��Ҙ�B���u��K6�iL��J�h̏�����b>]ls_�^3���kydVUP9����G,��`��{�/���}�"���nY0����E��C���;ڇ�ҊŒÁ�ߺ��p����-�
��SWUJ�����������Pd�rPoP�U���x۴ퟔЇ�H`�R�'�R��,g.��J�*Z�2|��L�����p��ݚ��D�+h�vZ;y�c)�`�O�A�Z��N�����fm��(�Ν�kT�A�����q�q�U��h���g���L��qI��T��X��_lj&8LB��w��� 'pG;6���~i|nWLh�9- �f�.�{<Nă�_�Ѧ��R�Q��?hP���U'��n���ʟ�n���o��zϧ�Pf���>k���G�S�� )7�������թ���I�5N��@xe��8�t��#R����',�D�H�	ȡDZ��Bj��.�L��E��O�B0����.g���%�niǈ�i#��.�2W��F���x\m\CJlCi]"�f> �f*Mt�sAF^#V.C�����բޏ��0^4d�)=l�څe�+;�H�PW쫽����ܡs-b�Sn$���踄��c�F;�iH��@>~��(���l���ऒؚzJl��2�I}�ӱзcԖ��S��S���-*�6A�Z��w
Fb��G"1�^��AE�20�*O�u�����x$���>�8�i�U��p�ͼ��2�]�ʫ�7���d�0�ƅ�RW���Wg�^# ��V�ɴ��uX�Q9�7]fF�55@ =��.x�|� �j�l**D� ��Ku��4�8P;���	J�S^U>+
��Z�*��KΞ;J����f�sEs����̜)w ݛ�[f�h���/���S�g�h1\��-����K"�X:)Nlo��r��1���~,Z�@c�I�g<�4���%6-.6��@�y�8"&n�s{,������I���UBG�r�ٷ� ]�����������:�I�}磊6;��'Y�2!�g��
������鿐B�������1p9 ���"����4�ȟ>�<�9VD�'������r?,~�l[�����p͘���6!J�;���n�}�t�$�JZ��I�G�����<^l��e��S\E~nMP�ٝ齗��q��$$���h�X�R����6��8�����hB�Ws�t%���P����|z���\E�؄�n�@&c{�[�9@�G�:�;�P��B�Ӧ��T{.*�g\��.��P5j6���X�Qt��A�wx�h瓭IPmY��*H/�+,zG���6�a�(f 1�m��ޣj�X���#?�\�_�n�ٙEL�5���
�@��٘���u���(�zWG
8��2u@G�:�ⶴ#Y�!ytbO�e�L 	��,�m�&M�Ps���Y\��?�9��J��-֭ Z֧��8��M�aKݟ/}} �s�;Rc+k/���+�7��$�8ӿ�U	�0w�I�jM6��Xp"�4m��h�O���O�	AC���d���?n:�����f/�{�$}_�͋�~0IWft�)�v���;�l�f�A�C�N�)����XMW^��W�O�&��,&�c#��f~���F@���֢ѾN��jw�[K�u��YA#ޗ �Y ��P&ữ�D����%x:�}�lPD|v�O�r�-W��̕?
��ix@ffR��vwt��4a���+^���l��ΰ��e~��a�œ�J�a٨=�:`}ۑ8L<�H<�t/GUu��8�r�����؝����C�<���S2���.QU�炌�����I������B�V�O4�͹U	��!9w��.�|_�'�,�K � ��9}[��	;�p�F*��"z��U������~O��I{��g综˧�i���?ۣ��� �`ړ���s�tg�㤥�tB /��W�l��V�=�sg���c��6���4n;k�l�j`�#�<�~#pӲq;1���RAH�5�
(���jg�5��̵�/1��
i��<3:�11�\�}���S�Ϸ�OL5�xޠ^O���)5u�R黮3Ъh4qzD!l�:FZ��=����W��ҿ�& g9��뭪��!�j��+�^bo3�b��������)���E݄0(ݤz@
Y5#��hjR�\�7�c�1�1�ΰ����8/�8�˅��d^@�p������c�e�̾�dn�k1P�������,OU�7��UD��U����@ im[���B�6�7o \1�
�z�D-]�5����x�Dc�Ċσ-�����˅�����$�'{Iٔ�����ŏM�Q
��np<��FռU�r�����>�/�M��׃��-��].����	p�7���:;��4ޚЃ��k��>���ʓf�z�<;'�܂��_�ŏ
�ppր0�����z�B	b��p!�?�^��(�+9���Z�S0���j'���U���B�l-ST���H��D�q�����t��^c?O�#н5� 2q����jJ�%���F��%+�:W��#�8[���ύ-�����m]?Ђ�1�����X���S���sw���Z<�E)�A+������`��[���n�u����^$���_�Td7���+ڔTT<�h��7@�^�%�z2�߮�_�O�1x��"�zxG�� �i䨧���ˡ��"�KO��]vh��nP��]����u�\\i��b�$�=�|�'0�����o3�E��1Ij)�[�_/��Gm�{��w���%/_5#���\�Dw�)������[A��ɉ�Ɏ>/װ�^u��a��eU�L����F��b���*��%���7�fo֐N�/���#���uΞANo��L�\^�}�%���1�I�z�c!=Bx�\4�5�.C���zL�1�A���f
3Ss9�G#�q��*�-?��N꽯Be��9�Oo�\+*Y ���
�1Jی��9���D7T���\���koG���食Iy�<5�/�5o�md�a>�q�ۓ���Vaf��E�Jϭ�P!9��S�u�|��b��7ܶ[�����z��
+)U8�kY:��	��|Y?�������H�B`�!4%"��ִX�{8�ĩd*"�K�x}����Y]%8�]��4�\2l�!^�����zO�Z��O���|�u#��	��C1h"Co2/m-��"�t@?uw��7��&?#���?CZ��\�*.W���Ns�'FMײ��C�7O�行���^�y�SЃ�f�$��ܖTma�]vc2+�"�3z��:��&&8�}�B�+�9- �����Ē_J�@��̩�J �`���k��ԣ:�t '�){x*����[[����n:��6!W��U'U��	7���43��7|��f�r�R�������8�'z�,�9�2D�� i,?��Ƹ����-��ၫ��W���Ӟ�{	�*!��H�V#=˺������0��;ț�A5o �EIU��3daj1���W	~{_�S��϶��b����K�XL�����M���ʄ1�k��@K'��"���_�09���}(y�6�T�r&��`�&���$S}�ïi�"�-�,��7?�?��<����2P�U5�ڽ̷ �&�%1��:�S]��F�ύ����8��#H@�;v
��Gԛ��W��7�$�c��,�=D���9�=ռ��2��ǒ��{�0~��6@:t~��I�jʳM������Ξ����Ls'v:e��]ûׅ�@��Ϻ$�O�zd��3D��]!��{E�B�!x��uޙAi�[9]�f� �vg�[@�ٞ�6܅1N)�<��sRĊ�P�R�����n���c~�[�ɕq�AS-,�G-L5�H�@:��L����"$�Q�	W�	@j'��-1��u����-�L��t&�5��P؅uy��1$? Dt*�1.��u�\�� �GV�P�S�)�+q�Gh�����[O�p�^bأ���-3�$'�ϗ�6ݵ����\f:1!�w�:����/�����"���`�m{�6��i�I�H���Ů�H�~��=�7�;����Tr���W��s֨7��������z���wG���Tr�}ɟi����}��U��-ɡEE 3�����(���S9x�&t)�Sfen��q��k-�L�� d'��=ë�yF��
W:ZX���vA�9v�X���ts�5��֡"^l�cx��ǫ�6�[����QfIpL�������N��k�ݚ@�e�eh�*��	�;c��c��dB>\nl�-9<�J��ul �:!v)��5>�By	q��_����)2���*$=J��eߕ�*��	�
,�O�r�a����e�Z��5)�i���Ԅ�om~Psh�T춋��V�D�D������6n����������E"�R��X@)�@�ņ+��3āܫnE��ݹ�W��`�)����y�r���a�HV*Td�%��1�ų���/��͉]�K��p���.�ޏ�����G��\�{�rnnMS��ۂY���#�MLU�qrp;� ��@m�1���Z��)�Ej��4`��Bϙ��N�_�'6b1�
b�`VC7/��4�$uu����m<�g�+��8��Jy�C�o�H����c����#�~k �*&��rh"=0��g���;��(�绎�&AX�bLd[��ڦ%�X��R�{�4�q�HzU5[4��ԫ	�|�-�{���:���:���wG�D*�R'ў���ոC��z��N�C��i���oƘI|�I��9�!���ms�P��pP6��f@�)�p��9�N׹^҉8nZm��Q�br�̒�.EF[��&Cr:��3��אM�Z!�b���9�D^�x�"P&Pc���]l��(Z���H-	Ă��ԏ��]��V$d�bq�j�xr�ʎO �`��Gnf:�"��X)DAX�B���s�����ǶW�K��V���p"���+_�tx_�;��K�/y� �	.�G��j�����2�,���Nw���!
$�_���X5�"��0[�L��G���@a�`�}5"M�ι8���5�|��.~�����t��93��2�E����V��I��k%'��ٌ]W5�B��Nl�I�sPE��Bn�V8��:��@���*��U��7ikʛ��15�g�cތG��ZW0����Z����z�-��K��e�+@�x����SèZ�:1߹? �C�q�XlxVHYEB    fa00    1630)>�ۘ(��x"!*5��>�Mr}b3�R�~��;
L#��>X��1���^��R �^0���,��[�%o��/Cz��@]'-ЯKTx��{2�D���0֥��R�ApJ�d�3���^���Ku��j�z>K��X.�>k/P���z�cm5g�!�	R�����)g1�<qj�7�m#cr��30L��"��-VE��@T(6��H��L���q�2L�e+d�_yz�ke�?hk��_�G����1����fyƛLĚ�]d��0��� �w�ba��|H
%��O��qJ�Cp�Yx5Q���}Bp����H�̷�^��A5�o�-BV �]����S_�cD�)\�/��V�W�[�=�4���4w6���{��	���©mC��P*=aq�L��ا�sV��G_XA�.��� �LzH�7}��ϟn�^��F��7�J?��c���� K�I|��&����c��=�Pe���%)�����ϤFY]�Y��;��>s��+��l]'nśeݡ۱�A��d����:�%����4���/%�Wt���T��\���D@7�"Ua�X0w,?����M�1O�A{o�ϕ��Mb>z.%]���:���$��i.��!�导�����o�Æ��[���5ҙ�{c���� |��|��H��m���g��
y�R5I�,����>o8�*�?b���ZY�P	�2�/�%��o��E����9sѫB�go}����<�����CA��w���.�xK��
x�������р�Ƭ���
	X���j�������=��f��vVrl��B�,?b0��q�4�Vת�t�>G��y���V�F]j#�D�(Me�~94�G�W�ou�
X@<�S����ƫ���>"�7BMK�%��>����a������x
�B( d�C#Ͻ5���*|P�s提�788ӡh�\�o1#����H���K�}@�SE��o�C��w����/�!�ܕsLh�^�����#�� �ABp�Z�ŀ7�����3��>�5��ͳ�O�6�g��y#M�m��S���hf�����Ǧ��e���KK���������s�
���G��ޣ&�ÎC�>�����v�'�th���tɔ������������׵XqjZG�-1����e�������Q2N?��cA��XV�x����U^��H�<��>�|�F7��<��(lT�3��m��M�q�bĸ,�g���A�����E�H_ࢠ�v��㗴��*F�S\>�P :��+�jI��xsڅ��؆N7P��Ѳ���j��H'S1��{�������`�[��L�j���J�v��\�9�܂=j	����*�q7�t7�ؿ �(��(�ʫ�R�\�����ˠ���zD���k�"�T ��W�x]1�����\�B����A��v��=�LH�B�؛�6�_��I��
q*���� �/�Ua{,!I���H�-Ge&������v��f�V�P3P�o4r;;wmq9��7��� CBw���| �MKy'��&���V�|Yj0��|�v����z����n�q�V^C1�k��O��!~�y��/��!+B��}��4�ǭktgX(=b�Ӓ5�ڀ+IzϓԿ]��i sL(�?T�zE���Ԭ>|'��W��V5t��F^g�/�|�����\�Bb��Q�z�f?$ac�;��r�y֒5�����ea��Lb���iC7 4�k�W����iZ%�����x�Bݥ�?xx��oapbG���,�u�Լ���sq�gL�R�p����k�[��lc=Av�ÎD�n��כ�}f�s�؋����i�-V"��>�J��Q��tN���������,W�/��y�[P[�m�_�$����J!!��_�SU��
�~���y,��� FJ���r~*'���K;��?X�z�?刭}hb�^Xp����),.| �Kb���� k��h�S��X��`�t�TҞj�Zpa9�u����S񁙹��`1���S��s?f�?��Zkh̹!x�[��������=�Į4^Z�	�7�V�6����Vm�k�6�{����T�}�ؒ�������U^&��-$B���ٺQ�U'�/�N:����ݵ���.XӋaz�Cļh/.�e���a���Z�@���mf��*�{��$и���U��q$�^��tn)P
��`˙o�=ǧ����k`�~��2��S�S�L��2Q��Mp���-�0o׷]�^t��++�Hl!dX�ʊc�Z#Dta?oW����;���6��.�Kp'>w�r_�}ל�g�5�#����5M�g9�*:��?���i��O{	C�QC�\����X�� S�O�=���Y�7g����|�9 9f*�XFHD�j̛I$�ؐ��C�]�'�*���H�e)���n%�$���&o�D����!�X3HSv�-���\o?�����J8�`>ۘ��ɍ�2���"{�p��N�%��V^�Ԃ��Pc�CxLG��P*`#u�uTD-��CU�]�ұ���z�N�͜4N��>z���V�P��h�*��\u������I�L�(����d�ma˩�����G�^�����,���V�[*���M7y�N�Tq�)U��&<�E��]O��1�WC�O7n�v�ݒ���S	n�٬�Q���0��'^;Ke���`%^��M���I�;��pɏ�f؍	59́�ݛ����
��=��D3���U ?%���(ܜ7�-�({?�Y�W�M��q�%����i�ګ�b�KAu�J�s$��Z�� �\���u�>���UV����vi�B�~1����H㼞�;}A
��2	�a�8�K�/�K��Qa�S���&O���b��\K��q�S�E�v^;�+ �u�]�/�e�v������b����Z�rޛ��8I�P�+B��T�Ӫ�.����������%דP����rYwV���Դ6t���.�3-���0�Z�{�G�"xZ����=V��j"!�*JX�s��40s��c���3��������F��i��͎�!$E�19#9NT�L��W�m
&jB.z��](ϭ�c�obǢ�,,@�.�L��!��;��(N�$����[ѵ&�[�w6���R���h�`�ӔpmF�K��Ж8;q֨����G~�o����b^�`v;FNd�L �#>��-�U�m��"���5G�r�G�V�a��V|��y�jO�p1H���B���-v���Q�E�!xu4���)Y�6�O{�+lF��-����i�^L���We� Z@Mpרt�2d�^@��-h��?�F���L�Ψ��1�=���� 1���(��5,��ПA4�q�P�+Z�Ƥ˞��Ty�'��	��#A�q����#��ز2Q<$;cqY���j�=�@+D�-��d~E�5
l)�
�o훎�J�
uπ�(Ɛ���Q4ټ��Y��6s�`����}��c�g��i�q�\�O�oΡuL���s�@@c�M��b�Y��I�Sv�W����3�^��+k��ޝ9��|	�v�o�+R 0���Y������@����<J�oC�,DRg����NM�r�o�����#klH엉+�:� #�Q�	��|8l�u���R#o?ن}���==��@��L��<�n�J�i8��HHX�����*��!Z>�e�\��L���\�5n���	��O��x7������7�;�!=�Ͱ���U�ӡ'dǔ/YJ@�J��C<I���6$)L�������g�4�p���;x��b�d���uOd������,bQY�D%�-)���2���P����J?ۃ�/�e�0)�dW����J4Nf'`�>� �_=�lB������
�w�r�&�_cS�2a"$��熜 E��1�8o�p�?��{sZ9b��d"�+i����.��E���(��B�Z������OcU�p�Y�&ټ�ӐG�����$�r[�i��0J���k�'��"=�h$��$�>���ĨG�Q�h��p$������'x���z����N��=dR�9�w����䥧�5_�2��C�Tغx!�u*>��Oê�K�跊o��Tf�DVq�aM��:�@�r��⎕bq�Gl4�ҋ�ʾ4$�|@޺�9m!8�����Q�}B�z�
f�/I�x1z��ܿB{�~�i��?����끲�F$��{��wW5��%v�0OEM��2��ڒ�!�G��]���#�I�&�SX}-�V;��r�s�J�c�A�b���A	L�J!o�>f��Ab�`�#�gc�[�[V��%%3�("�G�	4�x�3퀋���Ŧc��yZ ��Q�߰�V(��i��=79���@���{C�yMc�Y�S4:��l-G&��s7�sd0f��[�7�m�Rfz�>U3y;�j�ҫ
���"q���9�;_��E�2	<$��a#5$ƽ�O�$!�:����ps� ��:E�l���۩�m�Y�Ԯ���
{��%��i�:�ָ/��*Œ�Y�~&��/rV�C�q����� ����G������	���0�&NǤl'��V��u�V�~���pEm������-���+��\�x�/�݅�G-����w�V,*�ua�
�vB�w-o�G�h.�blJ���\�Ŝ5z�%���^�+M$��^j�LӃ����s" �S?HS�%�&�v�.�N��@����su��xU�C�ı�)7��E��C�3�2� �萮ņc�ߘ�OK-�W��s��Qi�#B���%�9�O�̯a�������4����	�H	��[��a�9�H�ͧ�Z��^H�-,�-��$}e�9�0�Ҳy'��i�JLW��BL����n�~���Qg������-#�K�:0�G,Xy���=�ya��TV�N�L��h�J@�ѱ��R��`�	��9�Vx�"k�kǖH2!��C �>n{�xK�EO�� Āh�ްq1�)�Pi���uQK,�/[�ko\_#9�b� �L�6ܖSR���Rd�f���2�+�fy���H>��m0�ק�Ƽ��y��F%9_vt^L�Ւ2�#Q%��WG��m:�����B�u�S���}#��O��P9Ł@�1�X��γ����X?�\�[�S2�k;ԡQ�ub���I�t\xD������Y�*�����5�J�u�B֊G.�=��X^���_���Pjq_Ԏ�W��D���JW��7�t�g�H�ZTD3Vy�N:Z�Ɇ�>c���G	�`9��TA����use�&G�?�p6�V��K�	��	,�P�dC�Nֽ��y�Lj��`�,��熳���Xb<%1.	����l��}a��^��. ���-�K�̫J��}���B����8\q]i(R�ec��,�1nE�wsW��>�6?4nv�}g0�����SZ]�x2C�)��a�c�����&( 	�6�آCډW���|�셛cZ/��p�^�✢���R��)&��O�`V�$8�>YY�ǔ�|��6p���.�*V\��v�B"ܩ����=<�to��A��_6����[���m�u����/m�-A��f�]�7XlxVHYEB    fa00    1620`������	�S[4�m���c=�X�"_4�E��i�8��_taXh&�������2�d$�7<����|E=p}�4�����W �>��׿='�"�|"���Sj�lM�U���u�گU�(o(a�Bc���jE ��xN��Ӟ$ǭժ�:��e ���KOK�q����
o��h�t�8�-��ϟND0�TPB�Q�C�m1(8�v��A::���I���l��pqO������Mb �$̊9z�ͧ���?q��� �����^?��&��Yu�{���8�T��h.�Q����$e��v�IN�����@�'���\x-�_�I���W�'���QS�?FI���拢(f��'?�8�8�~�����m���� ����,��n7P,tS?Zd��:�h���_�8Vk��M�(ˤ]��êM�^�g�!�����gz��K���ʑ^V���SU���9$ �'�y���
Hd�����S��p)��"�o�q m�6~ ���Z�:,?>	D�F�eN.v�N��F�ec���3-a�\Q�Q++���֡��α|ɩg�]�~����[%���2Ŕ���5�|��1����6e�65CBS���5g=/�q�����ױ�~)��y��Pu�>K����QF���7"���h\��k#O����O�Yf!�+Yȱ[ؚ~0�r����oJ�xvnkO�!�I��[�]E�%y����{��ֻ��ķ$B�,(�QSh2%��C���;K٧�D@k������r�>}�Q����O�t��:�ؽw\�B��l z#�!?�O9ՇYt�S+�ؠ7 t?s��7YJ�k�f�����S}��'���s:eL��B�)s.^�!��ڋ,��m�\)qu'
�wV:�؃��o����zP1ӄ@-8����I���|��*�+�P���IB	K�m@T���,@G�є��� $ M�-C���Ź׶����Dj���'L��S	�^���O`��	�Q�l�䳽����Q�>5�`nzoS%k^�ܻ���e�v��N(��e��"����%㢢
���N�/X�)�-��k��XW��Rц�=/]�
N:���6ud�{�Oǜ׵�kJ����ޛ���q��թ��0��"�Yڃ
��e�<l�kJ�5u����=��OP�m%[�r�X� 'Y�G~�u)��YUs�I�=�r�@	=v����Ē6P#-֜�j��!�WN�l,\3/��Z�1���s���l}�$̊�� '�8��S��j��%����?x^�(+�H�;�̻��_nB����G7�������n���}�-�)�[�> Ԋ!8��a���U�[�����]�:\�~-@���et�A�Q�5�t�CF��/� ћ^l$�O]��� ���(
i���SMꇡ{�t�;� �X�PG-2��&@-��z�����! o���}H0w��w��H����.O�}䳬�9� ,Ti�ׇ�%�,.����s���2N��.��bU�����d��R�' b�ۙ8T�K~�R��|�U7z<��RJ��ܝ����Qq]dl)^�5/�tk:��o�0Pƾ�9,GP���Z�vk�@8*: X���_B��?4�" ���������W��5�A����xYՇv���z� �X�7 L�U3�)E!/�(�i���� �.�*�"�{k�]Y ��o)|�����q��2��J�1���́���tE=k���_�/e���ly
������uÇ��"�.�4P%�j_���)�@# ;_��+}ް�5�8��N]:P��f�X}�7?23/�F��8w�����=� �����~�ͅN&�S̓��5"�3��/@�V�K��o� �Dt<�Oێkb�{��O�Qa�����ٛ)��P�@R���O�孟��g:�qMc�`Ȫ�罨��-H����7���j�Z:����Yt�I�HJBWLPA�"O�S�g�s���d3�U.��)lF�8�L��u��2C��j��W��R��I�T�P�iβi�PdJ�ũ�0���ɇ!O	R��P�.�h�9X�k$/*s�^Ͱ�>�c5q�����u��u%	�:��+|���!�'�����u�vX�Ɯ���L�~!X��j�(_HJph����\U���q�0��p���t�J�<��GJ��;5R���َ#}|�
�^x`<c9���`���oT�O�;���ZcK����7ދ����q�UD�t���E NU@��|���_1v�xN={�YdKd'�{�����PmƝ�0�o&�*�Jwu�i%��b���`- &���65��Y����z|*���ō��t�7��<���G\�ʏ@L�^�L!*��ӽ=����z�19�di�$6�	�fX��L�aƕ�0�c��Ҷ��b���X-��T��c�'"�e��d�� J/��A�f��q�Q�g�!���W����I�b ǎ�:D*�?�#��!�gH2�G6���a@��񈖩����N�BߩK�Tv1J��+��D;f�P����.]�T���ݱ�P]-r���F���V�5�˨hm#-_�"�,[�i�g�"o9m��(�F�iy�xdzQQ<�d�K���dQA���#�����]q�8�o�zW J�"N+R[*�dS+j��M��[ZfC����П����e@R����Ŭ�O���\��8/�j��� @��'f�@�s�$%E���,�=j�o|���j���hb����h	nB@vl�٢����f,��V���[ht�3I�8���7jyҨ�������i	j��� K?E:�#}���: �X��eB�Ҟ�Q{50�4�T�5���O�J���?���X�^l�F��r3{����K�w�z�����T3M=�M�
5��e�*�2��@&�z����y�S����	w�lM�H��C���7��׍�3f`�B�ʍ�Cp8�?:l��a��˼���Q�?�E~4�jюփk© ��W7��y��kX��g��e��PO�Z��ٞ��hN(��z_�а��s,l
y~T��UA�C���qL�T.��w��?Ơb�����ކ�I�>��ݨ��� ��u$�X��\#�YnpF�Tڅ����>ݨP����~�ې*ģ�]�a�1���sDO���}ߝ���/R o�>��ݓ��h� P��t7Q�0b�Rp���/)�ݗ���AW���hX9|C�\���ga4�l� D�$�U?���Ӓ&�?7\��i���Z��	��M�F0kt<����z����Kyx�د����1��"��
��X�~)N褔ęi3f�Zy��
�dhRbפ"�r���j��@6C>R6X��C��D�:��c8��;#��l|D.;��7Gf&���j��ѡ�jq�p����M��#�;�e��T�����\�Y���.t~��9P���.�Q.j�u,���=/X�Ј��<g)0nN��e�ޚ��tz���S
dWG%F'qK����^O���HC���o��e��f��囹p����c6�}.h��d4�Ă++D�hcC���nd�>��~fRc�݋�S�g'����B�?�8��	}UN>+��,+�]5�췇1�f�,&�S��'�L~P�.���Te�`��m�)�q������!�fq�	���U{c�; ��Qn�Rj�x�,k��`�S���=Ny~��-?S]�J99����k���E�2�зF)r-����)c�?��QaM��{ʏx}�| Q����Z�#d�7�Dh���5�Z	�dt���zp�an�%�B���ۆ�ջ.:��F�@z}��:~𫔃Z��d�P��{�R	����ܻj�:�\�*�P�U�srv4hx$mJs��"&Ŋ{	��!V�|�)B��X��ا+}�_#�CA���ط'(��9����I6��7�՛��<���ʒXH@��D'v��j�G	9�rǺ٢u(bO!�*��I [��a?O��q�\k���=d>��>�U 5)�Vd����g?m��A�����$�ه�`L�'��@G,������',~S�A,F�q��P����\Ui�����#Xx����l��k; �%�3f�$��X��a2=۠.}%�1G�m3 �shՑ�1�\����o$i<�����g��T���y/�)j��؃6�
oUWVr���o���G353���@�o:�%O������K���.��4�IS�\��{�����x<x (c
 ���:%�ɼ�d�RU�������Pq�v�S�b���9�����m�n�,81y>B�<X����&��|�V��Ũ��K���S���*���N�<0�j�-?b�nlK�F�=��V�%�ym^��>�<���+�sV��8C!&��QH=	FJ̼{�]F�JKb{�����y���&�d!�.$�fa,P%X�c���W~�D}nK��F2��*����t˞M��Z��/4Q���3qڢ���$5#MI�ttr{Ǳ=���}�k�s��$)�1f�$���������N�'�yZ>zu�u�����f�@��=y3��3u�Μ����\q:�
�@gB��
�%��3��8o��>�<�~���4�ؔ�`�؎z߰��$��InL!W`\O"�h�{��N&�a����lD凎�,�d���ط���_� F��<��7'��%"3�e�?�h�|��������]��8Z7f�PV~p,aϿ�.싄i7�b�j}�i���	�U��)�C��*��m�'t�>�=fZW��b�98��j�p2�dǤ����Ҡ��O���K�S�)���L˗d?2���T|���,k6)���U�<7�d��з�(���O���qAn`��V7/es̞�+��8o�`��)guG��Na�R�֩}��`W:��F'��S5[�/�h���&?4�hc:��`S�B���<a+ܨW��	���(�ǽ�CB���ȱ,��@�?���M���=D�Cv��m1=�送k��C���f3;z+<��·�X$A��f��ֱ4�9;x�=�-��+���ol����_l�`�R����
��E���Ҍe$�H�0	��B�d�R:�(�+��p<c���^�;���^h�x��zbH���iF��=ϊ��am�?��嶐��dP�d�kXl�"�RI�@=�;�Fųh{s�+�` ,Vg��?	�+��*�Ό���>�3�f.�L|�v�+��A8w�S´���THp�^n�羛`�щG!� ZD��/��'0�ˑ��D�?�>~��T�Q��_ ���&)�;ֈ�-9���6"����b�M��hC�ѵO�����K|9���m!=7D�Q�I8�^
�S�~X�u9��:P��X�f�H���b@:�*1�稓-�mcٕ"ټ-#���*�{38h�D��;1����A�'��1)�h��	����`ؓ��V�e).���L�G�0��f��kK�g����fG`��~�x�X'�՞�r���(�:�ʷ֜���
l� � �?B�l~���bΨn\���>�o �b�W�t�C��yJ�K/˓zXZj�F�D�0�t�c.)��J��j���_�G��C�ϩD��"F�|��I�<{XlxVHYEB    fa00    1630V���+<Ī��1+?_h��S=pvT*?No�3^"m����_ҳ��~[��:�ض�U�}+��I%?�Jx�&Y�1�36 <GDOѦT��2���xۖ�4�����Ky�V_��1�,�?�o�f�x�9&]r�J����u~q�c��#E>�é"�K��.�{������fn��E3҇�[��"]"Ȣ���.F!��C(/��[�6@V�4�����V���O-}Z�l�|���%����u��w��r�y�P�� Ԇ��̲�ϼ�X��!|���aO��zigp��_qa^G>?�\�a�mY���� ٶn��P��`�/�Q��D��t�B�_L�t��Q����ş���S��@�ґa���l'l�jU��e�(bTP����I�퐳��h��\�E~@�M�TAǂ�7��v5i�[�H�M$�	+-	h���G��V�cI-����?�\�A����\�,G=�W�-�=�@m�W���^���\>)d��6LV�+m3gQϱƗy9R�g|;�����@f�b��l)hz<?�!�:-n;����!pf��<��d�(@�	�"b�`5Ls�6�!.x;+p��WJj�`a�e���0Gg�p�,��Oɤ�?�,z������֪ΛN���&��e���0O��^.�6Ķ��� e@�ZĤL�	��qwբ��5fh3a>= ,�{>Qs}	�8ط!�~������������>��T�\����В���fк}e�z~��f���r����BV�'�?q�	�;]ߪ�7�M�6�5o}ST'�Z %Ҙ��'��3/��J�t�$a�x�Z�iʔ�.#���9 c�43���q����Ċ~�+p��锜�+I�%Xb��*��a{&ǔ,
Ǹyb�>2pry�C�렃��F�g�8y����$YНk�(g��O������/����ڒ:&���}{X�°�W.���5̈3G� �6E$�m�֣S�ȼ�"���^t9~��4Ҙ�Q�@���e�����$z1[����)dP���>�i+,B�ZJ��t�u�l�[�~gV8�T�<��W�;��~���73vE��l�G�v�!!���)$�m�~���z��R�V���FR��¼�$F/���x��<��[Ճ������҇ٿ�ǞVvC�y/D������=vմ�JC�t���l$P���ju����PjΠ��� �W\[���5�O[t��v��
6�U��2991��Y)57��K;��ػI�������N��� �ZM�Q�{.�6[v��D o�o���7§��e
Ade��;vߴ-E�-c=�A� �'>r�5���ܢV��i8.���a/!�*]�\��O(ƻ�F������/K�(�z�˧�p�+��~���G��C5���fp�o�-7F�$����-	���E��A{[���W��8����h�3���Y�Iz��<����ߌi���ξP+x\���r#��wAG��{W�h17ԗ�M� �����j܏���'���o�����6&�.4�f�Z�0bpӳ��CZ'�����O�J�:��3 �PF��=��/���H��9",*޼�*+���$��,	�O��ks�R<��&��je�� X��n��a%j���'Y�;�ѬJ}�����)1]�A��6��1�r�I?J/Okc	ɼ�]�eݨ�s�M�GR��6Y#��I:����l��'0="N'�\s/�������sp�hfMr��*J$�/s��~t����� 9���f��e�U�L�?2uy�L�GV�Z*o ~g侹z�W��u��~*�O�E.��gЙ��ib�u��j�@�(T�^������0w��"�4�j\s�`�~ɒ AҶ�.̆Q��_��!��16.��ck7lz�����Q�]�4��;�>�����reEJwN�,nF��fS![f��?2���sX���,�����+���{�������qa����C�A2�l��]��
��޹Cq��FS���$��L�D��JP'�;k6'	��[�C	"���V�=!x��}"nW�������9<(4�N�w[�����|��,[�=�h���,g�o�	������	���嶸L!U��+~WƉ�v&� �����68��)�@��ΆVlϏ�vR��U��p�b��M	�k���K���ȴf�L՗�?�=��e�������8�� �n�Gx�|����/��r�V,R��*�sӾ�k��Ѻ5����'DG���o�:�y~N`uA��sM���N_N50���&6w�
������	��Tk��!�,�	�j�s>[��B}�d�z�[M0P�=S��]_�ֺG&߁71�?v&�,[����߫A�XR$>���-e�>�x���L�Aj�d0��zU5���u���~�մćP�c>��8Ad?2R&��:T�^�P׼�y���հ��+?<��u�G��}��Q7�f	a�^�D�9?�W��a�æ��M��r��%B�%b;"��W,ʜ�	^�D�-��W{H�<v�U�Xǘ����_�Y�bI��X�d^��������K��A�|�H�:�]��)w�gcB1�!K���ú�G1.7�JT�FgW��_��"�N�����k�N\C��V�pR*�Sz�k�zJ������:=Y��D�C �wt_#��k�m5p��&��m�?/�)f	J������
(z����+��c�_�~�U�ăfק!$�Fx9�X�N$�J�п��#T�f(.~�@6ze{���{G�1 �W+�
�����J�|�2��7�� ��$��+i;�Yb%�i+s�FV�r�(��&~]l���9c D)�XD_M'�X����4�泦/�XW�>9=f3q_���=\9�| H;@�q�VM���i�z|��M&L�e�����
j����
C�o3��4C�/��=�	����:�lȌ=[#�m��fMf�'��<]���m�̯$��ƈ�j��LW�(z�<[�BM�JDl��vX^���m�"��0���<٤K�����V�fY׽�g�ZF�Y �xȼ`~=V�*e�48�k���:�(�L�lt�e��JT	Q�TY���D~�.L�T��A���W��B��l�� ������&�mԾ�èS�:dќ�fk���5��Ӝ��X�ɢ]	c"ǻ9VZA�'��W�b� �D�,^oG�]�����PW���j��^�$�X��9�C\O�\�)	��8pK�Go�m�_��Y�4�͟���sQ�X��+v�8L[|�|ʑ�ˤx�\�i\���R��e+Ѱ�ο��q�� �y�=E�
�9�2F���zԥ�6z� )�LP�>�v5�b��9��h�E�@u��k	7CYt<��o�K���\g�B$�SC	�$l�#��P�����ak
���{md>(K�j_�LT`�b�"�c�4Y�����e��3�����ԝ�4�û��Qw����!��Eq�quT~ۣ�|�蘸#Z~e��������� �пi
�G(<,/�۷0(���� �F�������0YJ�mbw.����iAB� �Ղ��P�F�t1�U�O3Y�P�D}*G3��ϻ��d��nC6��/��1�O�Ќn�
g�O��\�t�~��.���u�+v"�=����R�nd��T}�q��3'�ShX��K<�\��^�8.���Y;��y�)S�~�R ���I�.�4_!* �i�~�(9�+|�f����K)�(.�ر�l�D����PEܢۃ3^}��v��&��q/��E����*��Nw��x������}L��T�o�4����-��&ִ2��iEvwf�*�x�J*l�he�sB�_p;�U���������Y	8>D��Z�"h����(��'��q�ǔ8��)"�K0j�'�I$T�'ﱍ������W��;!�B<����*��5g���mm�T3w�l���ԇ"$e��\_�����6Zy�|��2��P*tN&v�5J=>���������ٿ�A��� �ݼ��"W��Rh�u�[%|�(G�x�W�U����Z���7�Lx]r�j�ٺ�`�A��V������}��w�����;����Z��eC:{��M��L,$R��A�ZЋ�u,�|�p2���ϤJ��2'>�I��|U�7��V���,�V���4}�Xn�٦nk�}��CH���N��
�#V��;��]_�
-D�O�Cv�>-��.����p5�f�ӵ�ogLe�2�G�����UI�sX��f�鍟0��ME�O撬Ɓ�ǺNV��w�5����TJ�I.�ئ7��)����
Tѵ�����Jk��$"?��33�� �y�I8���!��@��w�l"���'���MO,�Q�hFY�)8I�δYM��a�4�(�͞B�/M���2$�! �04��:�A�4�1���u�`����	|�[�`���U!�Љ���;F�T�W�ݰ7^H�LG�P]>��sA��p� &QT�9��[ᴗR�2z���q�2��>�:������Zc���馄�2��P����j<,R���"��Q�S">��ƋFa	T;�2׮��6��cvk��.���=������Ak�BUX���HF���k�d����tM��e{T띇�g��obh����<_D�@B'79��\��UQ���C�٦�.��sE�����ӂ%uGN� �s��Xa�<�k�>�.�����8hQ�H Y�l��y�ތ8�oq���AI���;HbA>ѢO�d���*���C��O��ĺ�2�����i�.%l
UE��[��� ��,��rvm܄��7G����=)'iQ�X��� 
rV(�G��]
���BU���k�8�W�B��Fyb����"�8//A}D���Z�V�OX.�#���-������̊�񮄏Qg�5�f���극����;���y=�_��X�]���I�i����ʺ[t��}l걩�i�d�z�i	��>mӻ�yz ��("������!67�%4�q�UU��#��:���j}+��mq�DĬN��
��$�7a[���U�2dVe�m������'.�(u I�@$7��cel���p�f-8�;𪎒�B,��uH��Y�WK��j^O̤��MW�#��MP8H�O!<�A�����j��8W��d��!E���������^�)F}!#����\(1֮�5Hj~��lR.��X����Į�V�E����Z��;���Eb Ķ�epa2���.���8й����(��'�m�s2��Dز�9[��-Z8T��C�y�c��[|��|���p=/���\3�����I` �S�q�#~\�ۧ=m����m��x4�L˿(G�F�Iu���<4�&.^�����VF����y,v�e���õP�`��Һ�'�Z���h������x@��^�FM	/$~41��x�� C��,�H9���O�v�JcT�`�q�Y|G���f�Qo���(��՘d?<��Y������z���W8U<!/�$i��q����ٕ뛖�Lj��Vz���»�^�D�;���?Պ��gh�p�����z}wm��4��8��х���*�z��p�il�.<:�:���_��-Z�r�9#�XlxVHYEB    5a90     850x�)���PU�O��^�\h<c�;�y`!M��к�J�NNXÄH#��Ջ�����?g��cT#���S���[��~Ei�3i�_=��8E4
)�d~�`*a���<��o*�@��!��U�k}+/�ʵxO�E�L@LKh����y�����GoR���$}+&�͈����v@@H`�Q	��T
��G]h��!��p��"n�Ⱥ��@x	����_ĘT+xFܠ��kK�IC�,����K�@�����2H+Z���n����ƪ��!��2�i�ȾO���0�h�/Ϝ,GV�G�H����ɡo�H(�}���ٗT^Kz!�eV6�s7�>��YgX�6(�I�e- Amr�4��ZJd����f���������S���6�[ên��m:��f�����}�#p���r��/�� 1������v��I���L��"��֪����_���R��dJ� �],;�b�����V
��@|d\���[�si18׻�7�R#��
v�� Q�ۑ��T�:{ �Ls���D�xbԳ;�z��5��Н=���d���AA�]�G/L?�����7�)����~�O�G&8���m��.��`*�T�5�'{f�<%V�@Z����S�h�{Bt����"��P_�m�s[j+;v*��2��;˚�lp�����5#���O̘��8֙3C|�к�=�Ӂ� ��@�C��w���K�8��YT*�&��ֿ�
��.�����h!miu9шX�f�Y��-�Ȱ"s]�.a����V�(e»�$�n�=HDCo��[�Ӥ�-��pfs1W~�p�Q2�Q������lI�k>�RQ������O`f��/6��`P������	\���A�j󤓞���	_ ����Q��f���5f�E,n��D<��UD����}f�b!R���*����"�^�&f�j[�_x%S�7c���j�s�-�P�-E�U�p��?�T^�i���W �ޠ+H}��s z�<*,A���-|(�VC�4�*�NF����f>Ҟ����ۆK���E��N���	E�H����Ϸ��J$���f�'5�ûq��M�nºl� �dp*�˴��"�����W��%�%}��q�ޏ��3Ѳ�̢�`������X��I@�.���'§�ڠU���O�W(hA���/�ׯ�̗-��E�;8%�d61c�������2Z��ʅ/*����Ǝ�`���0��b+o�^��3n�2E�q1�K�*uw���ېA�1	?~�4&�@����D__��4�&4�ȗL�N��s]=�
pve}������ݚ�K�"��a�i�
�x��y�Qk��RUָSD��C9�7#�T���[�=�H� ��2S��Yz*�n�b�`�#�"YD~�➨ڿȞ�IL��*Ӵd�斐�d�?���ݷ����[]�9�y:\��e̍Z��iԄ��(�q,�:�Q@;�󗵋!���P�������Fae�V���u�r�x�/U�//���Р�L�&a�0�'}r��x ��)9�u�f���u4��2�a���V��פ��/:f��+%v���IND�y���hڸ������O��ʮB�A�O�<	=�0�9��J�@���1x��/x�6�a2��3���x�����2ѳG�Y)�	go�s��JdLY4��Fϲ猣�Z�1G9\t��+l��&E*�UKn�&��>d�}�!MRþ\�4B�5�Ph�B�+M�FSQLlJjh2|�n\kh�� 
BdT�͛���06cg��~�EE?+c5Mqb�4�� TZ[����}����'��J"��-���/4Q�A�t,�6,�|f)q���'��E��������w#��kTLe�=�S#�=��Xz����'rGp<�Z�E��FT�_޸;�s�Q
6�=���`_�?^�'��\?KI��h�D@3Q<�Q������>�-�蕮('���U���G���C��iG�$��fz�J+x�>��Z��&�f����w�w��T'ڇ�ܯ��q���*��)o��?�,C�L�H�HYщv��S>��^��U�