XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��"R���w<�H�f�'+�"�31w��І(V�crV����Ɖ��#Al�ΰ(,iP�jAgό����	1�\C�c�%�Q�0�,Ћ�_0q�V��`���ڗ�i�cJd`��4(R���蔲#�yX� ����'.��1􅜔;}�Ԍ�#�؋��N1r�T����-�r�mQ��Gf�(ǵy��g,�������.}�P�cECV"4;���Lܓ�:�F3x����ɷ��oׯ�<�������Ɛi�Lm������̛�t\��{\�Qi6��� $H�E�	+�Z���|�;� ��Ï��&�D�K*F��DR�
��G��p�g{J���>iR�̝��x�^	c(�]�qM3�s0�/<�l���Ҫ��c��
PJ�S��c�,{o�p�P�xbSɖѽpLSrD�3�xbm��-��o;Q���>˽{'J2ȮŚC��M�_��x_">�tUq�L��l�̓�� �=W���o��>����"��5�}�)$K���o6�?�_�D�Y2�؉����b�0c�J�1y�>�(`����/���?�r�W�2?AЇ��W�T
9����p佻Ha�ډ�C}�������[�� ;'hF��߱ǔ�,ag�!6LDY!l�%������VB�	����{�%��6|�3+�lA8��6��5��L�:F����Ac�펉f��ͫ�g�S��Z	A�<Ȱ}�N�"�������x�߬<Om��n��U�J�" �b{4'bbXlxVHYEB    1c48     560Q��Xb�`q�"�C]	4=���h�qS��3��j�
��e#F�ft��G`C�f�m)�GV�ux�|����ɩ�[E���x�++X��_g�}u竡����,�� ��a:+�IejD���w7�(�0��u��"��_dAF�F��7|5�d~�����J������$��/��<��VIb+��	�p1����*���/�zH�\���UeAM�U3��A�d��F�9W��́�m#x�C�m�N~8��N�b�����2%�9���P�.����W��i�՟mm����%
�TR�dg�7>�1��k�T��(g�R��b].;,��+˶G�"�HU!�q�u�t�%�I"� m���\C�PAt�~�yߺ�֫A̐@\��M��N����,YЌ~��L_�YS��E���ܴ����yT��19y̲%��lR[i��[ɛ��*|c�Xˌ��E�͵��j�
 �;qj���&�'��U3}�}�:��B����G$}j3L�`��=_@�AܖuD�x�,l����߃3sf���������'߇y���R�!�m8���"�9�6~�9B����~�
Y�B��<M1r���D�<բ]��W
�d��E	#7(~d�z7m�q6Gq����q/��w8�����j6��f���0t2�dZӒ�'N���w��'�W�DA(n���-QK��6�R��
c�! R�'_py=F��=̚9|MӹH���4y+��WV,.b>@�0'N�e���rr�x���6R�'P�N�X61���숤==���E��+�}�6k�l�L��"X����X�,b��|unO���a�t��Q�z��ws ]_�l���>7*Ȋ!T�g����O��V�v9����Je�h�}w%۹?]%G�D`YF�`��-�Y�R�!���Dh���D��v�~����
击ZH�η��Gmlh�'Y&����!a�i����RՓO n�h��{C
b
,�,��}�N}��;�N���`��� �͞5X_X�M� CO</�`���'_�prn5�h$�6���Q�j�D������՗qt����v|\�����d��8ϑ���z�5Aos�t�K�@=�7uz5;tf�ʇ�]*�`���-^U�H�Y}��������I����BDf9~�jxӀ���ۤ�8��]]%���;���'9�{��B��S���
7{����O���:cq"&���0�D��� ؃*Ģ�A=P�v{��=Iye@V�̄�N��˕�!��f��v'��YNΛ���Y��F� ���yz�����R�3�qc4#X�]� ��^+�r[Q!y�p%k�rxs �[��