XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��a��!|����R�
_�Ag6Z����a5*��f�X��������3���P@13*E��X�*��ǵ\
�Ɯ� ��Q>ďL��2q\&XYT=����p�&��`�鬱c <fHOv�&���Z�p�����2��#�U�F\n����
	d��T��gQ�=�R�J�o�k��4ZP�p��
d��^B�|��WU�K���2��c����y�� _�&���J[��v�ebN��-�5�~i+��UZȐ�8(���/�yq�O�<5��(#J�:�)��5ncmrh�inB��7$t}4z��m���H�&8k{ׇ}�E_���0���F�����oːZ,���Z��� 4���B�t�s�F|*�y �jǝo��qS��z����o�EY꤁)F+yAr�+�T\{��.��`��Bx���a�*�0��p��|���5�|�_����w�R��Z�v�FʰK��&�5ܣ�Iy[D�L�#�~%��vl�����\�I�LL����N*�d����.��}�j�p���mKkf�%F�Z�V�U��'}��V���W�m�D�c��*��� ��Z�V�+������s�����u�v�� �/	�C~�x��0���M���βK$� k�%Թ����7�B�f7�]-^n��Ä#������&${h�����6q��:¶/}���\6�+iB_�Lo�E����Z~z���'���߹Ю�4oS\|�F�&g�p877����sv���#�V�Tu��=EXlxVHYEB    5ff4    1040���O4����P�C��S�r�}�-7-*�����m���7d���Y�����P���q�E��>Jߚ[ѷ��`-k \�����hG�ݬU캙�)-��4R��l!$�ۄ~/*� [R�q̓����
��E2]{��:�-K�2q�;���rj����d�ͽ�\HGc]�.��Ź0�-�z�	�\K�wW�㄂�����p���1�-����GDx�6�'6��[Ͳy��JD���k������E���,ǐx��I �Ōy�*[��r����l�� �r����{7�wSa�Cy'�֧��3C��"��|H[w������u���
@E������V"����K�c y�9p�Jv��^�͢A���   ��KϺ�3md��T����si����3�k�2,�8\�TV8-�UK�/մC�G�����"}ȝ�pߌ��y�i/}	K�\Uͻ�3Q��+>�l���r�ш.�T��	jg����x�7ڴ>W%�@�+*���؏쯙����C�r%p���\��'$buU��[�^��$�Oz���z�ú�YԘ$������G���~� )>+�Ow� /{�6j���9�H���c8�����(T�]���������%x�J�}ĖE)`�R�Ef��=����[	�ά�|4t�����j� )�g
4t�X�y�m�%$�����=:|6 �,�)ſ`��N)��OC��keҵ?G)�r;��8kN��
��N3��0:/o0����V��{�\I$&_�Qg��+��VTDr|)4���ӯi�:D*��Yu�4R�%�u��p��θ�1���[4?}ϔ{S��uk��8���7'^e�=�@��6,�~��e�X�#Q����L�Ru;G;FMr��6�7n)sB�3��#:�#��R�5!+����-y=��#h����9�,%U����L˭�S���s�L����X���vC?�����]��.�/;}f�w�o�|h�e�@3DM�v�	�����.���>H�^��e� ��F�>�۟�l�t��0����V���0ܛt8p57҄�Jſ��K�L�/ٔz�T�.��%)x�n����j}�	��lǄ���ʢ�kSw��u�j�X�����K��]���d�n�*'"��UN��T����X4_*�,�v�]l\p��riK��ʦ���͹VŘ�m�͕DMni+|^Е�������%��sYF�?��-�l�]�J���#]5ͪ���)����yp#R���Cn�pP���\rDP�Ѩl��63�s��ܮ~Xa�ܲ�}R'6vh�#���뚔q�,\�Ɇ�lH!�����}ߎ����*�aeGw�B ��֎/6��t͔�
ٶ��#�Ȏ���ֶ�赿^�L�6��Y���x�y����7��q62@�@4����}(��}0&	��Aj���������!.�O�}x3�_��ʋ��u���u�y�f�X�o~w`9QA�y�L�I�wQ�Yo�ԋC&<ܐ�좨��o���OP]T#��D�!_#q>�8���Y�dV�����zD+Ol~0�*��K��Y���%��N��K��tY�����c�i������ip^�7{Fx�/�+����pCAwF���?�ptQ��
�N������6��^���o�Ò��3X�n`&��Ͻ�1��(�^�"xj��o ���EL���ˤ-���N�5��ҥ}���	�Oѭ3�,NI�6TB8�.l�� ޶�����!Fc���8I˱�м��O��?���K4���鍊������P^���f{xV������ͅ��̠��Gb�"�D�-;3p��w�����9����-?���D��;{��0nOͥN�i$o������]���`��ki�x�����կM_�1M��DI�`���!�~RX
�`:SH-*3���8�����v���A�q|h�=up	�w{js�6��ۣ�+�I@��<$ ;��T��K{M3Ю�D;\(	� �Lp��TF��D_	��c��tx٪z�$%lcY�Ę�.g��rʠ�MB�k,s'�.�Nu�����6��*�,�	��Z�h��)X�z��s�a��5����;9��0���� ����(��i�Z&W���Q���E���lrёC�bה��s� ��GE��<��������,~KA(:=�X�䭺Lr�l	��|?�|�MJ>����3�#'��	�����U�����.����7��Fy����z���Z�W�b<��"	kQ�d/���ޒ��z��Cx�ɰ�2N@l�ܦY�f������\�_7�Hԯ�b����^m�:v	1�e���Lϒh��t�+Ǹ h�����xi�0dKY�(���/�-����ʉt�G؞r�B;��%��DR�̙��.!�6�DRfY�h3�`�	��?;��S��O7B�"\e;Y�C!�>���p��D�y��Gʙ���R�[$bS�� ��7���H�����e9�K�ǳt�`�#q�A��Y������2h�Ny?_糧�/�Sj��k�]x�jFeuE�9D]���*ʻ��IX b����=k�,��tpm4�｠�@zW]���zW�M=�Y�Y���:ǈ7�E�+!��(��zAI,c� ��
d؞���g4�[�	ä�`NB5���H]��g�K�,k��䑟�˔�A=���$d.���hL)�^n�)�v+,7_�M�b?5��*ʅљ틼���rD�`�́8S��b����3��2�������oG�b��[N�C��"�~#��C�����ɒ���3��)�l�F���䧼Mn5�3�m@u[�`���Z>�2T�|��\�M�"�FVjc����,�����A}�����L5 t)؍��n��cNV������P8��K�X��2k�*�o���P�r_s�\������Oв�w��cL��B�j��y#f��{k�O���C�0@L,����~ӕo'S�c���>�R��{����m�[k{�(���~-i��l���g=&�&��5�U��Xeq�KT�T��#��%`A3M��� dL�G�bC��痊s/v/Yi��<���yAw�QSu$U�ް�(��o('��ĻGI�PSH�ĀSN�����o�*Ѣ=�p�5�,��A���hF��0���o�,zu�Y��ut�C��:Slѯ�?	:fěߡ�W�E!�� ����)����A��_ o�L���%,�d�(�,�6�0����Tλ�׆�3p��|B��FQ;u����|XX3��k�C*;2��t�Io9��ևߢ����A{k�!毉H�г�3���<��JU�stn���eK	7Vה�ї�h_a<�kWE�~"7uW"���md&�Ϸ����C=�t,u.��G�"68%_p����l��%ITJ�&�r�}���u?&�oC�\�a[��56��Yyz�>� N�0d����@tG:Ed�o����eH�,�L~.A��o�6�?�uK� ���!6q�~�2>�8ל�%P/��:�K���N0S�Oon|.�NQ�h�7���N�F�+hP���?�[tstVN�
rޭ�q��'fD"��A��D+bԷ9O.���`^�R�w\=�����I�=�K3�y4Z��SF�Z���:X�P�H+cpД/�������E�<ڶ��U�-b�幈������h��3��}�FX���9����������IK?|���%C�Ofwp4E	4���?,��hI��w�fs�Dk����1�G�4���n(�8@/܂4u�Fo�f�M0�{��;�o�J�ky8�-�����ʠ�
�߶���{}g� ��O�\N��72��X��J*UL0X*��*�W�fΧ��c�^�S��h�V�d��ִ�(�2�������8�h(��.�4e0A�P��$4�ȏ� [-���ɉE�~b����#�[��!��5����^���/�P�4pU��Qp	�@/hCv4u���Z:ي��#���OE-<DI9^��팯��Pv�7+���1n���<�ެ�a�#b[��0E.!�I�Fr(eda��ٱ3�&u�Jk]^J|�3[=& �=��>�lֺ1R�M���u7t�a��9psdL���v5_��71($ؾM0f����F;�'<����؎����0kO��Z>��