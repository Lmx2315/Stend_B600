XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��	�X+�o|�>LM��k���%n�
��U������ߒؤ��O���Wj��8~�m� ���8�5kH;$~?�g�\!�z[̞�N��[v�jmw�Z���
��;��L��auvxJg��o�?|��!«����Iq�iyRZ���[8��%[�z6�R����=¡>��+��	�)r_��E!E���bn닅���g6�%��	g�dg�fe�[����s��Io�뛞�[�F%�q�ߒ0<��1p����k�;������QE����zrF��}|+V�B�MŜ�g���q��k:�؇i��.���{�ep��A{I� ֎��ި����0���U�������&�	�8�Ӗ�g�1�'o:3t��J!�����[wRW���(t?��#x��<ɾ��+9M��X��*��˹�;_��n{�V��	�hCWh�4����[Y/�us��.m˗���+q皖p��??�;2�����J
f1G7N"m&�!̥t��{��rHU1�-Г,���x �%�^H�W����	��L�Y�������]�a,ckY�G�w0�7����eV�	w���\�xiJfu��lO���Q�����Fo���}aD4����LD�rNW��5'�񨊃Rؕ̀kj�.���k
O�R�M���cwH;��E��$��-��������C~> ��w�[k�9�@���h&�M?�p&����We$��kwn	�!*���ep���bx����"N	�c�-����\�s����]XlxVHYEB    1d4f     7b04���Ռ8/��5U����&�ٿ�}AV���?�~��͒ۼ%��.^�Yk�պ� v }��,����ܡ���#�񹻒E?3�.w]�h����4���h˦툑�5,�����]��<B�\�ۖ�8�f���g_z-F�΢tZ���u_�t�5��]z��Pj��\]���a���y�%��A]�)=a$��<��ah	���#�!������jӍշQ� c�3 ho9�p���[Ϯ��(-q�R��Ah��\��8=���x��!ÿ�=n]��w�E&��p
B�����[Y�������T)�����'!]� �W�f��zxy��HU0f�ms��Ð�?�c�B�u�[������ir�؂������E��YK��VM@��xs���1����]>��������r�GwZՌ���t�l��y 4S=�s>W�iu4�L�~����O4���q�-���'eaUS�+�e���nA��<�J�˼��q�"�X�wV�����B~y}JR�ʲ�*k�y���.׆k.\t�[���*5�����H�F5�c(��и?W� ((�ZT�\�eӤ�]�+X�Ev���ٍ�c��2{w��9G������1U��#�.YCܯ*�N����M����m�+�g���| ��w)��2�W1���#[^�|4&�i�k���F48Q���0�|�����~�O�(�;��
�K��mۭ��y�~���{J��qQ8䯡�"l�|�Y�~��6xY Z�n�'�͗�c� ��]a�")U��4� �H(��]s3��ݬ{pp�Xg-%i���@�)Պ��`ïK[��9,&g�>
P��Ak�ө��A�jM��{ֲ��d�iԭ��1m��J>ڈ�@�^�͋�2�M���屵�O��9���G�b�yN6�CD�Zu,�Eq�ƺ���@b��{���.��!���;����P�Y�x�$mX�V����1sv)9J���Ȏ�䬩"Sə������p,�J��Ŵʯ�f�5�J̫$�>�7�)3�ai��e.���M1����y�^w�jQ3�(�+,�|����A�h��U�k�{�*����|��HOD	��hh~>�s)�붐��˖��9f
�&���C81f�l8{�����H��"L>�/$X���� �')�E�Y�7~�?���|"�~��=UA�.N�`��v��3F#��꣝6,�~�l7��[���@��![�U���mÓ¸��Q7�`CmcL	���#�g��x�M��@y��$ݑ���tS���f��F���rub�9ԇ���ׯ�6�X;���g�	�2O�C�p���~�3��́�\��X�O��7-Ħ���ɸ�D�Ks��p�̈́��-�J����=j=d!�e3��+��t�kU��N�U �߷�k��;�Y�g+�P�8��eO6}�w���t�N8���vU\�T=*�r\#�{K��G:5��UZY��� ���<�f��g0�E�>�toq�W��1I|����r�/lVX�0�o��A�_��Taƥ�����<K�����I7@�Mx�S�X9Dq��M`M�8d�^�э��|w�7��X��:�=�,'�y�*o�,a���]���$��-�i|�.W����?��_��z5��\֝I,)�^�L���#��EyBo�vS�B�zo2]�ެϞ�6��ڠp3���1�+L�0�]5���?T9t܄uN�v�(�"��V2l����D��4e�[��e�ۛ&�=���u����,��@���s�p�3���+G��ެ��AY65�d�����e*L���+������y0P��n��e������2����uMs��T�U>��n2���)�oND����O#��":i�a ԫ&{X����u�����;g���w<t���'�7�Zf��P9h:��3�s|��O� ��I�V�I�R�BI