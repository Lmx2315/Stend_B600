XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��W�����E��6��y+l$鏣Ic!��O>v�|�Q��O}o���M�s��	4�<�����sCT�?�w��<wO�(��l����b�fL�;ݦ��h�9�
�/��9�g6����)����~��G��3%Di��c����=��pB'��l�h�Rϐ%��p�?������6���9��v͉�7I��+��4�?�Ҹ-��l�z���f{�Jm�'�r�h��1��[�Ob�Z��
���Ҥހ�@�1a;��j!�c�&���j��X��'M0O �v�p��B����*�[;)��x�H��i�HE��V�[0�SE.�]~,w�P/��"�oҰ�'�c:na��Ab���9�ָw���Dw3��Y��rԪ�E��M�U�|�W�C��7c�����ü����U/�&b�,3[3��ϝ������
ioI�(禝�<���^݉���������B:i�qh�����P��y?��`=��%`�Au_ז�l� Yh����g�v�$����}�{gx
Y\���#aFñ� ��N�Vr&oe_�K�I�q�p���q k)��p8��$��cy(w�x�H�͐0jg��>���Vdz��J�K�yl�hl�U`�vˠ�LpZ�#էS�%(�Ԍ���L��r?���g�$3�^��?Bz��J�.)n���%���eP���/{g3k�#`ܧ+����n�d�mN�ۓ��PrF�N-�}��=j�x���X����H�� \XlxVHYEB     7e5     330/22���r�\˫&L���:%�!\C�c;l�k��ސ~�C��zJ�x����K�b��nU
P'�R:=�������c0�wbTv����y�P)�:?�åOZ�+�xn�@߀1���ω�T]�D�y�����拻�(�U����T��+��BR�0���ջFT��A�߃����x��9Xg�C��i�5ˉP]�Í�V�:�5[����U���׽��T�NZ�0Ԫx���Yla}\�n�8�XtT?)v,�̆��5J����+}�^���qQ5�|��._uIS�ż.'�K�}>���Xz�vA���ZvO�hn��μD^nBP���@��)��}��N��P��$ҟ�g48 ]/�z(%X�l����9��!A��xTDL�`E�FZ#7ǡ��u|�7�tO�x�'�3c�ߩ�GS�w@�'^�ED��8�����`@��)��<^u	�� ��O�!�\�-�w`�{v�G�ߨ�q���9��9:e��6�����(q���lQI�`��Ğ8����}/��7�#I����Yk �K��ٓ���6�exl=�6�.���?w�e���f�d�,���e�^��!���l���ɮ���5���Wk�û�)�x��̟Xl��Ft��6����{�<*��' bڨ��6�e�$;�5eq||,�5��=�(+�GO��*�>*���'�Vy�]֊=抂�C���I�W��j1��p�&S`�|���"�����Ǎ{�ב��eFX�
$	j�(��G��C��ٲ�m�F��+��-��[�u�C�[�N���Nk�o��RA��C�6���b�^�d��