XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��@v����+�(�T����R�ܪv��!�<���>�i���;�0nt0a���T(��M�=,�$]e��T���>��/&����bΧ�Lq\Y�m���y�8uA�b�˪iO�ҷ#P��I�K!I9�C��Æ\�����p���_�=4
^LlsZF�E#��$!�σ��*���y`�&�hO�>:\A<�7�ݴ8K=���3�x�FG]��Cϵ�8
�u�0��v�®�(6��m���\�)*�ͣ�B��'��A�]Cv���PE��*܁{n���O"m��@ᴨ�<hΛ� �ek�җv�*�Gt��@�a�=�04�4~�T�V�������=�ք�`ǎ�;�Ⅻp�@���~���>�v����Vz��ͮLR��QMYw.]��|��\���pEɃX�Qq1�r<�~�!�mF��Y�}�K�V��q��y��,NcIqA�O��u��)��I"�[.Q2�U�4�s�TP�`Ѿ%��Y1I_�{�7=Qv����"T�d�9ꕒz	��GC:�-J��L֜=������Yfy�!���v��t���ަq���ޱ>ړr�������d+_�_��<��7O�K��U�y(({�%��O)_�j��P0[�7�Q�ߐ� ���	q�~9l=��@����9�W�r)�D�tۥM���J����k�	�-]���\Kq����L�v��F[��#ᑟ�H7�����eF� ��E>�;�u��]�u���Q�V:g0I�.Y6"9!���֧�o��XlxVHYEB    15c3     780;Qj���s;s�T~�q:��"T�z��`S��b��ոisW�y֔���?h�l�%��y(	�<�د�c%�q��f�U�����a-+n��ĵP4k���9&b�`�5m���'A]��EN�_8�%�`I�u�2���D�_����S��}�f\n�z>�谹~I�2I|��m�=.��;,�����p($r ~�uu$3����%����-!t^4��
joH�-�(�Ml@Ղ+�?@q�#��-שּׂ��������Y_�<�Q]�|�q�qѵ�M�q��[�]Oҡ���ۨs�Jn�����Ɨ�a���X��v�靸��?���&��^�G$�(�x�Ugy��ǉ�.rԙ��۰�&7�V؝?�
=���5cT �jE}��ȠP��\�4,>����B�p��u	:}��:�!����[�.^�����Z]d��K�x���=_��T ˊ%�+�QV�N�V/&�CFHC��;�xK�c���@0\&fp�5��9�1�A��c���k-5��j��nHnr�n�)Vp���(^�%`�Av�� �A���,rY��y�7����e�il�x��n��{���y�����)l��+��3x$��^L :='(-��%3M0Z;<�%����Ƅ�%���s���F�
E#,U�� ,NG*�F4*��l� ��*���B,���4�)�/?����N4�����$\���)�ğ%�!rry��ؒ@�Y�ρ�A?�*Z�,��A00>���
e��^�GW=6�����C`���[|���-�������e�%�swcn�4��C�-�fS%��&�&���z�@��2%%��u�"������奈�zo��:�Q XO�PR�����K�ʺ�=l|s���D	"4�P.:#�B����Ŧ��StMMC�����o�xC�ؠ�W-�+��,�/A8 ��sKv�����W�ʍ���0��:D��.`��b��k�G�"^�� ��=,"h�^A��S�л�Q�ѹ�� A����ɠ�݂���[JI�&�Β�Ԇst-�I=֟<��U�6�Dъz*��~��l�T�D�{%#��$[ޯ��Y�jv�ܼ��[�s�m9�Y�������^�T��ن��󁘰j�D�0��N�9��9����/��Wsm�W���f�{��Ke_B���rJ��@K��`����/ݣ�U�����H%�N�7���~�]����)@�@Y����<PT�nrߴF`O�>��oo��Ek�̞��i�U)|�
��@U����̂��>�i {�$?����\�?����#8���ֳ�[d�*C%g� ���>�Gb���b�$o��E��I\�ip2���Ey_ؒ�<t6K��s�镮�����8!%��a���zY�j/�ctdaM��ץ�%����5TG@���pd�wm+笅{���lD�[��^C;��DeXf���HE,8�B�} .6uJ5��Ҥ4Ѓ0�P�?����%��t{��n'f+]�$�yB��ȝd�y	f����ZT4��;��YgƬ��(���!X��5N�_�+k�1�6P�%���ō���O�Y���ˬ�L�~D�{��#h�	RD}�����3r��U M�lj4�1��J1]Ā�ܚ�&ċ���9�ޑ����h��%x	�/��s��D��_24 �k�V�����
�p3�� �3I;a�_�1��@>�П�=[�+�Yݭ:4�_�#7�?ߺ��5��I�|0m�(���_��!K��Oh t���'��~��bh���oP�-�?��S��T�ű�D-c�i[I%trU}8>�׿D!Z����+;_����p�.	ơ�8o��i]��f��V(�x���nػ���W@������k$v�~�
��]i~D��/w�ƯВ��B\�]� Nf