XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���.��Ⱦ�7����OUTMÃu"�(��C������#�;�=�}��׫i����mr	~�)��hn���'���R?o��h|8�~&&ъZ]�?ɦ_�K��l�Ů^�b[O�R�U?�V~y6Bܯ8�X�/�B�@���:؍^Hc���H�k�����=��X�}�ս{=�B�9����3-.�FBk2���2xL��o6bl�2&��<�����>7Hx��2 K59'�(O,u����zm>��D����U�9�ԩ���;�&��K�$('���ߴ%\9�Eâ����o��i�3w���>����H�)�}|��3���"�b$��ճW���#�se�m����UEON�dZ��'q�_C�x����&Y$�g{��e�]p�d8��4�b��1Pd|��mlW�I��%>�j�5�w�#/wU=i~[�)W{�}��K?'��eO��7(�I�=$�mY#�]�e�DaS���Pη����<XE���h�f��mܶ�7�8maVD,ܥ�@� �%��"4_]o�	�"�!�U��s�@�������w5�i@L��N� ����qx����O�����l�g��z���8"�1�9�2��E���&���5	;=��l�>k��n��0
�2,W|Ob�+!�u)�tps��$ݏ۝��a��C���\HX���!tH�G��!�����L�� �����Q$<LzC���,=��*�K��Tv����R���AXlxVHYEB    41c2     c40�-��� O1��.B݅��+��\�_��v+�i���0a��񘫬��@���\ٞ���LQ�)�����g��k��B��E�p�)j��c �G�7���p�����4����<���ip+r���f�}/բg�5K��7Jv�])����h��ƱJ{P��%ѝe��vv[o['��|Hwe����0��m��pHT�O�/�QA �o���EV���G0s��FgEA��@��/[Fq��-��+�9�q����1�Fx~��-M�I݁�Z;͊Ol'�A���y&r����w�`��7p��}��_��4��Q�6�j�(�`=%�<�0LN=��#W��ӟg�C�����YT�PI���M#�5�^�% ���Ԟ���М��θ�����1�woL1�=��W�,�e{�)Q
|�ې��êx���&�cC@q�$u+�1%���\[�p�������1d����82j�}Ɋ  �H3ޕ!�t��Y��mz�{0�8-���V�n�̪�$��+p5⪘���@|(�6K��>
��u~�@uYR����;��f�V��H '���vʨ���$C
�!.�U<�\�Ui7Q��A��������!�OI/T��NFԚ��S_�U�n��*�bþD�&7-$F��	l��l��(|kɊw��'���M�0��L=R�����dtPFF�aq���4Z���z��)��-���b���]����WV���6D��P��� S����S�=���*�LLs��V�!����0�*����Z�ތ0��"�z�8ag�"%d�P�8s���*�*�zf����9�Q1?�tЁ��ZI�C�<g��x�=��������$ǒ��2��ZlDc#b����@�� 	���yۇ>�¡��Fc}����{읁���0����!�æ�w�B��a�}4�uSk�����s+7��� ��L�!��-�� Y���yIݦ�9�c��h������7Z�k&����0,���@��6	�p�C1�}�����0�U��3�������lBJ�����K��An��3P�1��Бj���"]C�3P�۰2���_��z���o�e(L0^4��8����2U��r��SYpR*��U�= °0�Cl#׬�!��<	M{�<�ԇ �/���~5��}N������86ʸ3c��C.6��?��ۃ��,�*+�ŏ���N�Z�����d��-�$������#Z�gM�F��X�u8��T��3����x��tg��Y�1�	5`s�k��qJ�u�e9������DL?@Q�g1�qS��}���d`�޷$�H1�j��,�d��c�*3�{�_�"�+�ݡ+�޻a�^�;�_�v�@��6�������v�5ƚ����|�~�5����4���J�բ�k���K/F�t!Xt:A�Xc���
�%��b�8�u��suXO�MY!2�Lc�cBMRB|Ht�Dc(d0��?$l�)I�g�_�0�B�������>{�x��_�@by>&`��{fs������)����h�n9MB�{ a	�y�J�9y[y	�a�6���	\&�h
-�~����PA�`;*.�h*���EW5�r9�b����^ ��2�t�I5o���j�V[`p�9LT��o>޲�\�B���E�t},ʵ%С���+F'�D3x����N�NP��U�#�v6�~�1�'���fj^s��H�S޳	��9�)\���	Ly=���yy�-ՉwRC��\�(؜�ګ{h�̓.
h���Lm��`J�/�Q���	1W����鉫��A4�p	�L�G�_��������Ȭ�ȱ::Quɜv�����	9P��z
���b*�~5@�7J�N����5���
��?�(U�a�Ͼ��(�-�g�4���F�<G�C�l������~(��\u?������]��vS�nPp���J���mf!�t�^ �L<vH.�LS�O�#�-����Lx$-:m�ɵ�1|�pٿ�|���t,ö���3K�o����U<R�b�W�ԚJ��"ʺ���@�"� x/�W�Rc�?����cD�ڪ������QH_rD-�Ɔ��%�g J���`�d��JX��zYj���J�������2S�(1yԈ��#%��&TLe���w�W
ĵ��<r���y�r��tV.�b�~��=���
Lyj&�U����@&ի���Vxe�!��H(/�s�u�ꚹ:�����.FTQl������ё9���2�H��Ϋ��k4��]��
hdo����7���}�v�<dzB�kj��{2��f�@�e*�/k���_����n�l�ɄJ��!�p����,�Q	NW��q���ԯ�`�3b�]vf#{���a �'��,�h�&^M+���iYgF*�������aZ�+��\H�����D���M�wXu�VK���FB�֊���0����ۏe�/@��i�������p�D)������W�&뜢C���xT*��Iȫ%�t�*y��,U�����7l�_W"�=%�c4���Q�}NF�ɛ�Y�/�[�,�	��qz�iэ�'����u��cI��YU4���	���!�E�+��؆P\K�����U,i��?8�]r&��P��3��Nc���R��	e��������N`&2�<3����}sqX�?�N�h��ó���(��Jd��J�����ОP*��Z�m��$��
��q�Q�AR������!UQ&�ly91{���ʅVƖdw�7�(?�o��	x=�j��'^~ᬖ�l��I^��d���z�2�&�Y�;?�'&�2f�(���8�P`$'�
r�� �4I�(Ҩ�Wr�
U�YIݸO>N���Ғ6kI�uM��캛�G��
�s ����/}�U�>ॻV�r9��3����So��d�t89ϒTT닟q���ֻ^zX��U��6��˶5R��m�Ҳ� �\Z�sx,�_4�;O��Ƥ�7U���&�q��,�^�.Rš�&�ь[�SVQqtQ�������VJ�魰N�hSp>���l 5	]u;�[�WV��O���ۯ0dAv�S�)t���t�7q�'�g���<�������|�މ�