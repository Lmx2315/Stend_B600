XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���7O��O�Iz|�s������e2e/��ǁN����Q2��P��Xz
�0��z*������h%s���6��]�*��S*H��P�e����?u2gH�[��=�U0ID;�l&����@�	�$��)�U�̃M�L������Ym|��ͤүi{F���������WY��S+ף� (��n?�g�<��ӻԖ$d�3��1��f�1�L�D�,���1`��h��!U"C�m�WU�n�ɳ�fc!O�f�*��� f�~ͅ�-�Н5���,z?��h�ݙ�Q" >O��$�7��H�a���y�61�
��i��L�|.9M����/y��w-�%�p2��G�qb,!g���P�Q�wi!���xZ*�D2��{?�F��K,t@b�p�0C��
��S�
��6n�
T���x+yDr9s-��oe�i��S��_i4���6�?d'��&q#�?��icF��v� J���H8�-N2�g<�5����z:F�Q�|2��68 C�Y��@��o"��\��C��y�1cRo�ׂ�S�8�%�.��l���_�@S�EƳoq�q I�u%
:��93I�;+{����U�mf:<9�I�<��Tf����F�������� ��G,��g1?s� xt9�VV��޿W�8��S�hs�Y�R�3,ʲGD2�G	���3�ė.�>��`�ٶ�ƗAX{ٲ3M�-(˻lK��~"���u+ 6�R&����Q�b�����$�D�E���XlxVHYEB     7d5     300�����cư \oG�g����DP�5��`we��Cj1PF=�� 2r�Gq�	��M?�ω�����z(��/����
���JI��p�)�4A�#<�k����2.�����ed�HQ�r%�{�2i-i�(�V3/<N��������S���~Z���͔3�=.�O]%˄ 0��FB�S}QXQ�%]�S���I~���()4��	Y���������;Q��RAǅ[}Y=��_��qґG�ʒ��a�f�(.�+�Hh���.B &�v��K�+�p/(��WL�N�紂������&$�(�H0甛�#%L� ��3\�[�Ck-����Yu�C.0�d��ⶦ�|o�@1NJ"+�'\�������zR�:`Z�Z2G��ɪ���Z� ��[�oN�# =c|y!!A;�TgO��T�`�M�~����������y7N���i/��̈I$�9㖃�jS]�*���6N���q�]��%����0p�Q��gni�����v���x�r���yb�����A�:���'/�,|B�$�z1�趪
m?O���G�eu�$_ix�m�ĕQ��t����G�	@����[��6q�)���?�0c�������4M��A�<
,ڈ\�����v�~i�8jU�O/�[�j���aƚ0خ�Js6�Xa�P7�[*�է�@����g�\&��^�f��l�o�J�}� 3"��AM�����K�%_�=��i95�7��m��}�� �[��7�MG�g- "�m�@�ȵ�4�����