XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Гۙ\h�,6?�B�y��ud���;�k.�<32˸����� ,�9�--:WrT*�j�Xϓ�����@��'(��g

�:�A>�Q�T&�f�r�� >�679a-�7�QU�γ���:{��|��嚭y�)�2(��j���4��FO�z.�V�;k���ذpb ����i�h^��`��	�1��Ey��'�1 �����&��/~��U�o�uD2&��	h#�ͥ�U%�v�QT�{H�e��B|����v��zp�������]8��[ }x�����x��aZ�!��lv�L{1����H'!B���P��^�A��yo?�X\��
՟�sl��&�6b�_%Ϳ��^��h!�T�uU�r���>���i��n��b6�S�d�?R� �6��L�\ b�n��H�z3��(�y���d���1S�d����t�G�9�S;�C�o���[� V���~��eH��-�2�,��5�����:�n��?sGt9�=�(Я��1#A�I��l}�غ���w�}�1L6��o|0��
�� !�+���E�o�#�Z�����a��Be?/��~�W���Z���E��JJ�����6ưY��j������^(�z�r���$&Ń=�*)��u���$X3j����:������,}nĘ�V�ܷV{p�C��12�"LZ��qlZdn;�J�M}�̸��T�*34��h@�޽���}�I����y緷�3������g�L%���DY��~^m���XlxVHYEB    3c92     900�[�\�HCz��po�1��ͱ�m?Vù8 ��k���˅�4�-��K�f��'~	L�J��>|��n[���I���A0�bt��������dihۍ��X,��Q���"���{�G���R���o�
I'��8|O����0���q���\�J���^�u���1ۍ����ߓ�W�jB��W���b�	y���a͵>������_���.�ziĵ�`%Y*��
u/� )���p���uP�Y!O���V��>�k~n��a�N�J��BY�bMha�Z�ހgv��9WЄ��;��Q�]1� #��m�Rc�H~�n�W>�
�	0B� �������Z�S��q�/B|�7����ϲ�XV-���S��n=��@w����;�T�ޟy0�W��%.Ώ� X�P��;�{5�.�7���5�|�p�?d�IP=�E�^Se<Re�z$�mz�=js��%^�fhŬ����neV���ﺃ����YHk��\����qe�E�=w0s�8�&�jmԆ����~?5���S���!a���	����	� ۃ�d*C�~�I����P�X/�έ���|��t�3~5i�y6��`�Ӏ�	��J��_�|0�4�=Z���Ř�d?pv�����,��8<!�t�3�չ�Wa�e\c��_?��:i�r�M���i��*�k@!+@^�KVh�t�I�`�٨@�a�)�z~
ԓ�*�8n�>�l&�Fr��&�J�! 3kLn����r�dg7��m����U�h�C~��|����~����q��`����N0�q����E�g�V��>��G�ˤdzu+S�y�/��S�`$�x�7(����%�����P��3��dw2��;Y����/�J���C
5�.��3T������ER,��F�����T�1�衳��
��U��S>K{��3I);�6���Vc������D*��1�C?���n09��%�<�# 7���o�C�<� �ֵ;ey(��Nl����-I<n�U*F_�2J^����j��3��lA�d�8��n?�5��ܙs���j�&D�F�;H� �e)�xaF�V�d�¦����md�h�$��x�a��*�D���js��-��:�4����I֩��>�5^�̔�JV���7��BD��ܨe�ͳ�A�8D��Z��	�u.�	JW��=�B��@Wm+�
�F��Ί�s_eP���S�UCVb;1i�B���9��F}Q��'"d:���#?��8��nQ������	[�}�@�VPT�1	�עt��)����2f1��.5�2h�{�W"�������$\����
D2�˷�7�����` +=�ٟ,��f�������RQj��|���7��G�]�V��R���Q��D�iաb,��K
�D+[X�2x^���B��)}g�L��'���
�����f�����|ǌo���Ӕ�����V/�6'x���~�wk�11�S�9��ަm�o�N���t�)N����|<�[�է�[����v���%��u��L��S (
	�a�=5E( ��8mB��pN���Zn|��_ly2HE�qH�R�r��Hj���x��fx�F%VX�Ԩ����}��M�R�4��u��o�Y�y��QNEȋ��d��Rӥ�Z��ձ+�9�������_ ��@P�Yʹb�I��^@�/:�c3�����a���/
VsZ$�E M
��@�����O��\5h)Ì��`�a��}�A�t�Ϣ ���M,Nsh��_�<G�.&��ڏr�� 4�*shB��r)�b�gI�K�� "SN9��!��gA�\�E����O�:�U<���H����G�	���'o��( [ ��K�|NI.�z�3T����'��17l��+����X/O�<b�9�|ǀ˅x]�,���ު�{a��\s@v��Gfǣ���B�yNx<�s3�m��x,�;�N�0.����mXg��\��EI��.�n��[�ω5Ͼn��6��p���W��f��K�[*���	��ߎ@�0$�5�pࡷ���ϕx5��EC�I�A~=բ>c��}0"<�E�
�TY�e��e�Wk�$�;�Ly"��D�\��2�|7�#��]��&޻ɿ5���W�I$��88���L��+�xӨ����W O8�T�T����w[�t�*)b���'���xg
4�B�(n֍�_*2����"x��Ư�*��@l���r�b�"cF�62�Ҧ>��`�6	��si2	���