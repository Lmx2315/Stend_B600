XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��5�k����:�>��x�L�3�iB����pƘ�{�E�?����hh�d*[)tT�v���i��s��q8��Qi��Ʌz9V���1�#�[�"�"~��x��f�x���|e-!���+G��U>�LɎ���r���~��v���rt���N9�����`v�uWnj�^1[�g��i"��"����D�wurD��0g�жڄ���;T��TG��B̄=��Rk�WqA���<f�n���/W^�b���M�&�-i��78�k�����B����`@۪l��B3$"��o�{b�x���(��B�@���ʳ�
�҂.!�n�6�#~`t�9�R1�*ۅ�xꕿ������s�K�?(�)8%�JX6N����eo�aI���k(۶󜗾�˭�������<�l�d�dEM��D�4�(��G^"�X�<�4�X���J�HCiEƐ�r7G���Bx���Xx�L�z�zweS΁�2��r$��$ٜ�𯲊P�4Gķa�\-T�?Ƨ�gk�hA� ��8�3垍'��CC:�k+���3���觼�u�!mD��y�'\�
y>pO\���J>�2ҌoJ���� �ۂ���Y�F����ז6��Y yk��VY�#�
�+#�UC\���T��#���fôo��uq �Wf�oWl�/����D{�?>��2Υﺺ}Z�t���<��W�,�%���x�r��W:ҪwuvD8P
Ї�� �,c�g�;��#^��[�3;XlxVHYEB    3a1b     d40�OjR�#��h��'�*����b���;��d�p-*`��ȥ�Xo���歽j�aC̈ �u��i��� �j��1뮞a ���z`V���� �<-:}�c����l��]6C���4k��y���r��/���&r�6k9�_*��2x��l,���Y�~|2A!�N�MN��[T������e�6TNZ��˪��Lj�=������:�];%�ձB��m�E�i\*7���)2&�>�/��:�PtV��b&���b�_&"��OaPG˫���%�z�i	���l,B�������nY��݅UJ.2\�V.�a��� H����c�R��p�2��p˝V�s�ͦ����:y\���3��#�%@ ���Y�I������Xz��Ka��׸A��ݢs�٘�T۶f_'��������e����}��MCcG�����L��b%#��\I^(��\�=G�l�ޮ���Dtޙ�����q���cL}~S��FT]�j�y�ê�ܕ<T�;����up�}�f�m�d��N-��}WgY�}��-'�N�Cw���!��h=��$5-nq����ۉ8*��0�|9�c�K���u_���  �&�ko+�0F��G�q=�����Y���%��}�E����[m��yD���O� �T�����x
Ѥv��S<X����8��7M���w��a�9���H�]��o��{�$n�R��Z��V[��s��H�	|b�E	�"��	Њ��ݰSn>����� �k�νRLi	��A jX�js
Y�Z=8K54r���Xf��z/e�*d���C���cr�x�ti�\���4z��l�+����Gl7�NS��t\���#㨎�����I#i�Q$��[y���}��٦��n[����{���x�@`���7,�ݕ��`�\��y�w�`G�5\��-ݖ{BV쪿/�2�MW�Y�A8�fM[;_��q�J	�'x�c��y3�eZ����9
���0`G�U~���S(��w�a�DF�7�6��x#�c4P�
�@�M\�9��+��W�s0�M���{�����(A�ҷ6���ko�{1<4W�����g	(fI̷	�T�a�5��Ў���`/hS�2DR�v��fr)G��h�'"Ui'wã����i9i�?�7�X�FNN���v�r?�]vf/��.X`�{5�L���Yj�����p��)��苸!Oi��Șe$ ���8_��ȶ��#��ƾۿ��&+B\�����O���0M�bV�3�~��/�;��&r �~�sz�GoNcМ�,�a��/�@�e�;>+"]�tî!RZ�d�� �)ud��4d��d8~��
`��`w�܌{��Y���a�����T�%��72�������AҊ#�Ԧ�h��ew_RneȨ��r@^��P��0�����]������H���*�g���Wo-J�4�R��K�2Z:��U(�N��-��Bs�<KFm���4Z8d��f���Ɇ�u$#�kq�p3����6�~ݯ���w��������-҂R���V��j�Dk6�-
T�}.�0�cp�tpK�u�)N~��`X����a��;Q�rL{�Ve��~�d���x|bZSGw��#���j;�QѼ����BW��|�P:�|���,N������M@Z0s�9p�fiI�|NΧ8&9f���]�N�Yv��"�Q�@��RU�Hz��A�j�� $��G�� ���B�+�;Nb!�I��v�� 	�j%�����N�l�Vu��"�#Z9��U�����b0��2��a�:֍�8�����s^��[oq}�&a�|��?�f�>=��U�"�K*g�#�@�o�8�%����F�a{/�ܾj��
�^̫J+`&���s�룿�b�\#�l������M5���	�����2���s�&3��y���U��š�,pPyD��?Q�M����8�3�D��j� S�x�k�yfb���#�x4�!~ �<m���N���m��X���L��[�Iw�<8.�S��"yw�T�빇JDd���^��o�I �Q�˒��c�gL�E���HP����oB�i�X��\���H҆u��;q���Ȟ��jrY�٭�}�	ȜW_��z3��ƹ5Io��0hW~�i�%p0
t�I-����|�#��	������3�4t2����o*@��N/--�]Aҧ� 0�#�g�4&��G�֓�����qr��S�����|���:��!Ղ�Gc�Q�N,o:�y46������]��5���h�xP!�L�#� m�1u�ml�6�����_T%�|NYL��|�v�F?w�Y�^Y��C�`��@�r�3u�jL�4�QFt��YU��Y���y�'�k�����kw �[�r�
�Ӭ�[g� ޣ�5���V`��<BA��2e�2Ȅ��2�|^)�|x����}�	x|�Zx���Bw��6�嘦�����J����'g�Rre޸�����z �b����*��t��)�;��ͤn�&Zc��PәJ�,��$��:{'n�����
x;��p�����Csw#���Ը2Sg79_gY�o�Ra�Qsٮ[�JR�D����Me��~��%��x1riD�_;[��*4A^.�!��k�1���^���9*\��i���M�g$7�����+x�DE�K��IZ��@��X�[HU�\���k���*= �I� CP�0)�>;o�Q!�7����Gh�gr�Y�/�X�����f<�\u���^m�*ȋ��vg�M��>w�+#o�b�2aH��!5W�p�+^���UY�1iO�����R�}�hy�PUS��N�_�qj2S�b9����
V@��޸���దo`�Z�����õ7M"H����@�t\�@����JaV0�stJ���7���X��B�T↯�6�^�!����KnM\rn1!���1W
4���1g�"������2�݌��g�6���o:I�X����jQn,�V}�Ԁ����/��3���������S��"�s����Ww���a�eHі�Nn��i[����~J}��t�,fXo��p"=�yA��O��]�=2H�pË��V�S���M�S3�CC5ȟ%qY6f�#���k����s<���uq���
LmG��~�ڴ�,���'����X�5H/�4�Wh�0$��bok����\��]��O�����R�x�|��*O��0����/����U�9QB�x4�T'yb��6m_�Nj)���<����_hC2�.mӅ7����¡��dr\[�)���d	��4b��դ��\_oi��۟��4����[A��j��h�������