XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��K5���@�P�D��w��(]N���-_a`��&������r3v�gy%B&����廚'1t���Y��Gn�ru�%Y�=-���Ay'���61� ����d�q���e0ٷo��ւ����t<�U3�ґ��J�2����Q#��cx����^�y7�!^.9O��ЭQnџڡ VB�$�pŒpd���������Y�T�c���0�?x��
���=���8�\}�������t(4���<����F|{hL� 6q����e�����N����O��)_|�~�E}��<j,O�����>��p�4�jSk%���l�/��:"� �R�(V�c�p�� +����]e���� Uq����=3O���j���;ct�ʎR��.��ӿG]f�C����]O&���{�U"a�g3Q��8,���5�o���'�,{+�������Aܔ�nZ�Y_�p�w��=�ćׁ��ʞ��hK�g1
�oZ��;a�PILCvxI���rk�>��lԿ��/(���r�Z#�@��La,'D�R�t����7�QY ��>Cl��>8� �J�����o�vG��>��u�	��aH�,#��R@N��o��+����E��>�M�;=	EIi
�y�'#3��Xl�y`*�z�)�D�.=999�;�Y$^>3�(!*��"^d��v�4K���.r�&"�eq����9$���4��I�xD��x���8e��b�M��p�1X�%���8���o��ttGlQ���At�q��(?XlxVHYEB    1f8a     780^�����1�fӠ |P����(��������ܹ�ʄA���qН��X�
A����!����w[ڥ�xԋĞK���d[T������.��~y$r�H<��B0&����3����g)���7��?�`Z.�('���nwʡ.`��W_�ξ{��d�6�j����C���|]E2�+7��Yj�Q}cd�=p d�!����yq���'���([J��@6�3�����e��4!����_G�PT��'�"���6� �v{U���\ ��p�ϓr��w�@T�3$����xj:_��z@s5���0��{�v�R�s�=<t�H�X��^V�|)��$���&���	�lu��Bw��~Z �)r���	���Bl�Ҵ��+Aq%��~���w<z%~^�`�vsV���5h,���I^m�"^4#�:��&��A�i#A�����g���܍I�&�M�i���i'A��$\4;��_�Ww}E����h��8��z�y����"�A�1p�( �K�ZR�l9�NM�\�� --it'm��8J��l�p9���܃�y��2�K��YxtM doiՂ�&��(c���c��L���������I��:������9]�S�_}�����Lw���H۠�>sf��P3��˥������رy�B��S,\3g&����s�����.Ns��Qx�>�J*�鞿9��O���K���p�` ���::`�S��'�f��Ղ�
��~�
Vi~��@ٰ�
nX_m�>e�0P���Z���K]p�}��B7N�%�
�,��q1
�A��P�SQ{0�7�9>����)T#��F\��6}*��+��sOs�mH��8_B��Es��:,�߈jq:8u�JS�����#[�����DA�*�}�O� ��L����� g���U&��<� �-���/E��'���h��W��Q�4fR�;Ҝ;�YXo$�2?�ۇU����o.�k�3�=��0L}4�v�{͇�[eO ��4~�u����M��{�P���ׅ=��B.}+���H;�甤�P�/Ў�S�|�咉���Bf|y+^ۆ.�GO�kK����l7�@W�%/"��=� ���.�閎ŷLFa�pP��|ep�҅:�1�Q-p�%Ȣ��c����L�#��뙴�V�m�h����g��X�-���cl��,�����Xi���=���Ζ%��w0��b˥S<�@ת���K��Gh����՗�'l:�W�7���Ĺ��>2I�g�f,�L�
��ҡ	G�b�:~�ye@5Hy�a���������0c��xp�^�FyC/��g.�xR'���q����p6���H!�����&�t�S#��n5S6�0)ӄ�/Ff@�����ә83֬����V��jM�9�8J_0�c-�O�6�ƾWKϏz�������$�`q�6ǔ�&h��4M�]\���;2��df�����G)A�����Y�����L˨�(ג�v�qs��w�/u;w
���D2S�+,h�� ���6�v�^ǩ��)Fg���Y>��Svt���2�C�Ĭ��,�Q͊Y�@�F�m�|;�h��7!dU�`U�6�K�JYoy�,��Mju
���+E��9צ��M$k�P|��R��i�m{�wBO�{�N�g�mK̤Fk��E�v��2�i������o��U6����A]�
9��B�B��[B�x��O3�h�o�ٕ�(��V��2bn���_���u'�B^Hv	A�8q�%�~�8$?��b	ܟg(Me�N��nV�Y6���a UPl�L���_�I��Zܳ�i����$Y�l��"��͘�L�A?�ܓZ���%Χق[N���~m�o������ÿ	�����˒��I�+��o�J(՞AD��@	<���g������