XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��a>d�GU�Xd\��
�~�Dv�jmR�#U�U�EL�u�P0�%t]ϐ�S,�thJ}�^�K�r����$*�%�½����N;�1�4"Q��+S�$������f�#y���fB2���`��G���`n��ڇ�@3�bCv�$��X�.ϴ��p���\�O��s3c����>��z��t�]�/`L����DSs���W�5s����u�UT�vl�9�`��@���M�9t��F���.��Z�^�K����ˇ�w�j��Y?�y�(V�����A��.~/�x���k��O����p�bY�|]���I",����`:�C�i�˯d;>���iH��֏R���� z�؎L��Nܾfzq������ŀ��#NA�k�j3�{�V��0m��;9a��$J7W�3A��U��YhC�E�ʟu��b"R�ω���16�q$4�����ժ��^�ԧS��o���@Rc�1��j)�"�����.a��m�/���R=Zt�/��ڜ`L���+O��T�9"j���NPIM6S�o�D��8M݀:�)�I���{̵)���i`�S��o_�d����u=��}��s���XX�b(M��V��*؛��5u߄���)a�&�i	�o��,HV�����:�Z�႐�+`�ΩMC����Hw ��G�R�mQ,;�ȵ]d��A/Q�U�u�P}}��t���@Uwԅ�m7���;A�����I�zr}�xw=B����\�%N�#XlxVHYEB     705     250���l̼�4��*OW��'9-"���4iiS�#�:�����8̃���$�U��N0G�"&�]Nm�����}��/���6�)P��%a׽�S�Ǌ���ϡf�$ ���x%�r�&-2V�BY�a���o�D��PXU�cF�2�d�gu�dg��5�"[�k�0�~����&fHS�/�#mhX��PY�x#�9����Q,*'���Oȭ�^FR�%*�B���������R����2q6-p�D���x<g.Uغ7���ۮ��.��0���B`�	w��������T1��8��'[t��!��VG��0b�ڝ��ډ�y��+� �$��kO��m�5�<`��7�Q��{%�/5��/�T���ǃ���~���îy͊m���,�X�8�m:��gI,j�Vh���+�K	Laʄ���F�����*����"�-��7\R�F`���O�Ќv��+ͪ	&![��F`���:(��x���I�]��n��gK����jj�
<<
mx���Q�t��D�A����n���`AH�o���(�Y,�=��kZMJ���$bH�W�E�Oxh	�LQ*��8��h�