XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��I�y�1��BB#��ߍ�P�o�9}�`i�/�D3���_��;�����g���͙��V��)|�/�� S(@�[.{�sv�E]�NX%(K���#\
�3�R�Vهe� ��N����_��>�$
���,h�28]0w��~����[�AC�{����ݲ����ދ�iD�$?�螈��%�
 r2;��"v��؃}�o�>�f���~D">А����(�H9�����2��~LY6�����DsoX�.G�̏�x�Wp�"q�1f'�ػC��`
v�9LJ����{;��!{���dKOH�<��$~��Adr�,��|-�g�V�����c��	�]�lq�sS�M���!u_E�ШHW:-Xd�`�]�f���_������Zo�����q����1�i�H��4-,6SF�,"f��HT J�f*��運�`�b����5��}�8�+�T��)��հ�s�_C��I��'9�/�Su���|����#�� `�!? @hj�
��x���t�R]E�9��j��b�l�C�M���	WX(��	8��m�tc�m����>��D���L`����y���"�h�IC��@k��]�+�]�*ljA�`nu�ў�i��L ^��9�M�p����sܝ��i�VR5�)ֵ�4�����@�ٌ):[��P��3ٷС� k��߹��N7+�c��݁6���4�
�*������-�#�}�� �^+P
�v�?DH�}��8(��Z�:���e������|O+��k2h>K�XlxVHYEB     a7c     440y�+��êAX[��*�Z%�7�-�{_*��=NwB�β�|�TM `n忝I�{�8�wu���xsF�g�8���Լ:������?��P�'���d���<�x-�?�bF�`BC �F�
3�h�"�ȟ���v"r���/�_l� I��&Z3�:�`Y������hv#���/-�.��g'\5*��k�+���k�>	8Mٱ72���;:p�o��� Ǘ�X� �3?��D�`�!��2����v���ߌ.B�?�'k&XA;m<�@vaO{!�Q?2�t���ٌU��5�7�ogW����+���;�,X�>I�ݴ9,�~��\��N�<Wb��F^e�г�u�L�ulou��1c���a5����_iAS��R���SG����6�d�q;az
QC�$E��{��T自b> ��=¥pA����aAkA���G�$[���?��i�P!��P�UY�W>7�h��B� !�DeP�v_i
�UB`Si�-~��` ���\���m9��mɝM��W�7m@��C�h#��P`����I��i����3�d!S��Dlչ80)��;�	���tQ>��+�!���.���x&+�� ��#��X�}�F~?�/��2&t�j8��We�I��$�5��O[�iW��p����qh Q�+�s���b�i���e�eaX���'������a��͇-^�3��MX��鋆^D��D��y���L
�6[���Lkgr��Ao��o ��Ɓcp)U?ة����W+6��F�g0A�%���0l�68Л�d_��#na�h��թ[��R�{g�zYn�N���x9z�p�}�É��',�t D�3_.���-�szA�H��Jz�}��~�31��0a�������4k�1Όl�@Q,@��*���f׋��\�<���X�o��ܗ8w��ΗgːӚ���'�x����6����uvuAy���c�-DhR,8�[@N��'�<�s�b�Z���Vm�:�X�ehl�Q�;��v�u���ǝ����?X2gl��?o��:�*�Cph�ĵ�뽪֋��\�f�