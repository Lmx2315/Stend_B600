XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��2J���R˰AF�g�^�;��C�XS��Fw�}��C]�^���5��!�4B�VG "�ʉ��5��9�ؚ�UR��vQ���j0����8��fŢ��R"�ˠ�ɠ������JsXC�cy`�=��h��V<������p ��րJ��Y_�*+�����\:h5��⌉��_���K�����f@Ta�p��HOM���[�:�!���P�$J7]��#�0��N��EQT��d��S�{��������-em���fT��2���hkb�e�����'�J~w������z �xm���Gв#� O(�"=�4O?$j���h��{P�`�v���v��!��P9�B�gE�AД�_k�);x`���~��&A?i��7W��8y� �J�2;�5����k�:ٛq�F�*ʼu�9�`h�:>4�_�jD���������"��R�M�i�*D�雧��d��m�<�D�[�s��茌�#���S�#����d�[#�5���x	�p�0N�S����g�	3p���LZ��R��[�F�Rr(��'%Z�u���)��|bT�i�fRS��M�5�y#7z�/�N%n�U��w(�y�M�'�_@�_e �0��$���TU�y���ݐF-��=���&�4�o���V���w}5�bW�����7��O�����d잲������!T��/�IHǥ1?5�#0�_;��#��P�DV��	��>4yD���׹���>��e�3�.)6;����GU����:XlxVHYEB    9944     fd0�)��w�zN�c��%�)u{�怯���Z[73�<��T8ʦD?cdF�BA�L,�xl�`���5�V��0w����.�v�(x�í��m�c��쥾WP�:L�i-?� R/_��O�Q���o7^�
׌oK�I�w�C@�C��녌��(���*R��i4c��H~�~h�s*�>G�m N�;5�p����Q?�Y~�#�s��Lr�C��B���(T�A0�����5��_���� �OqZ#�~���s)�nn����i}8�-1�ᕄ�P�Z����꺚L%\��aӷ\�5 IQCCǼ.�I@���(O`��7�U��tz������
ѫ<��!lma�zg�Co�u�,*f57��[�/�3����I[d(Y?���%�ڥ�H��X�ZX8����hd%: ����;������O��#y�	�x3?�:�;Fp�zb�RR��C�tH��W>�=I����'E�`dz7jM��<��H1<����6�)���p�C@�����7Φ�S��8�?ܳ���_��n�駍K�aIA5��OU�P�44�����GE�T8i~nt�K-��Jqh�Ų�B���ێս
�X����-£�/Uu1��l��2�.�?ϟ*�)� w�_�KM�Y<�P?��GG�v+]K�y@=������	
��BQ*�T��-�Md�ߒ�y�v8�=�#���Ӏw�� m������d{1^X�?�rT3��
�K�t���
En\��u�󏮹L4� % tb����t��pJG�)��@"�u���.�l��2Cs�_�>-�R�ǜQ3�� �+]���S���P��:8<�Rt��4͆�WW�ɭ�� c:�]Մ@\�F�RYS%=�Z����K��"�r�?ͯ4f����<]��Y��[�!Ϡ��Ǉ@���o)AC�yw�����[�[u4 ��K� ��vQ+���31C����<�@zt��5:�&j9��>��ϥ	����r/��V36�{n�׍Z�V��%�z=ٸ��e��o'֥�̂���9�PY5����V�u��>�nߖx#Y���'"F	�,o]jp%dq&����+�㠜x׵��@I�`�Idv��I3�_�pZ�=���{�c석����¼:/��-UCإ'=xg{��b��aE�����~�F��y)��$r��[��}i;\ p@�Q8&�
���'FlE���⿚�1�s��Q�?x8�H,�vr�6�%��f<����>K�Y�p�����<$f�#�3=_��=����ѵ@��&�ih�l����G5\�R���2Kсe�
�Sr��ߓ���F )�_������D�T��FC8V����vk3)�3�L�$+�N������Z:"��2��8���>]��B=�� bLm�_�5�a4��b>������4V�:^lH7�Æh� ̠���<�u��Hs�⨿
�WtS�75/�#�9��ࡲ69H �j��tz�}R
�BO���oD�ލU�$��"!f�qF`�C�4�6�'��@��;L%�dՌ�P��\uu�V�" �h�L�(�K�L��<O���ب�^:D�߶�`�`"?��F�w�V7,�Y�j����NYl�x&Ym�ciU�AƚoV����J~,�xp-^	�q�NaC����8�QM�ri�B������n7c�m��������\\�8<o!w<{���׋ͳ<&�S�	�n"S�F���������,{#DB��^�ނ�o�ώχ�R}�kw�߷>|L���d?}2���x�a��5W��8�Cu����\1�32r��#Rv$F���[��]�Sb���`IT�ِ] ŊM2Wc)�Nޅ��|�	xnb؍�}cL��'.�%��"F��t��+0z\F;�O>&�>������Ѕ�%��꫏���`��O�C�/L�1!p�3z%>>1A���Y~�����Q�S���_r�3�Ռ�4U������1�uW���ۚx<�h��g�r�Zq�39�dS��u7�Ǥ���2�Th�+�u�}U��{O%:x���jM�9�u�����ݧ�]��	�8�q�p��Ä~خ�nCh4�Vj]q����Nn\�A6�9�0��>�9�bMl���]�7NH�^�e>��QU1�;�.�1��r���6ϾlM*^�_ypA�C?>�F:ȟ׬-u�^N�:��;�|Ӥ�����
b,_=�3�8~��j�t�*U6�1ErWZH��_�/p��tٙ�f�X00��`w~
-��(Z��Z?I1e�4�J�3xr16����G���j����4���x �"�=0��ZDb|J"�waf̢�._��U�]hw�ʉ�ok{]�W	J���Ox-��ĳ�W�����J�xhLx�;
^���{4��J��Y��h��&�ڳE`�:��V��X5�Pg�[e
�؏�a�5���,]ڕ�^��L��pA��	jݍb�,��>�c���8����ka��˶�V�_Yb��O#��O�3���X�6���!�IH�9�eg�x�Bo�J��`8����@�dH����E���ͧ�E���}R�R�7��v`�&��K�<U�2`����<��S2�� >?�7�H��:��M�ή�@?��w��n��2�$��Ϗ1}��v�W����a���%��(�6�Fh��ha����{��`[5�h{�|�E�y�I�h����@��6��0�7}?ˮ�ɵ�Y�cF��h@�>�/)�/����Π��.�T�w�b��ၽ@��F�F��k �'�����5�K��7���Z}j�fU�Q�˓�_��(Tm�UPR�
L��E5榛��s}��(�Q��cdtc���)[Y񂛖���m���~ hF��>�_�Q�w�&h�c�~z�sb�C�.��[�XY2k3�%w�Q��S�uŮ�����6�rx����ך>�'�l�R+R;2�\(!��޽�Y����;���^8J>�6V��=|t�Y�JJ-ܳ�m�j���/H��YZ�����������%�>��y_��CC����-����,4�G�Hzww�E�:T����0��S�J���I�Q���%���ly�s\�'�v�rQ��d1M}����臐��-�.�֜tn�?�q0�khR3vu~��w�H���9]��²iŝ3W�ɓ���=[\;6��g6%"��D��طx��O��!��E���g���T���=����|�@��w����k��J���j���n�nR���y����yCL��Ę����[p-���M���HQ�cQzhiz�ٖ�����]n�[�2����ܘ��ܟ��q�Ƽg~2�w�9���2c���MZ��`H�W[�n)�,XԂ�^��Ƈ洸���2�m��	��Mi�T~)чr���
�g��:Ye0��o�,�V�F�[�N��bk�ĝ(<l���M�19�����F��?�G#�<�a�
��pxX���'�\Z0s#�ZW�Bڡ��J[~j���+K�	�]��O0 ��R�`�����U6Lb��������e,�ZV��c�V�g\ǫ�|�y�1�R�,M܌�� ؝��G��~��qgiĂ��K{�w��5��*�aT�Q��Vu�v�q�[vW�(�����H��K�Y�⊡<�6z(�G��x� umt-��9i�y�IS6];���=����E3C�ձ�;�1�w�:��R�I!��C�H��b]ǧs�~�R@��;�S���x�}]��@[5D88�5���0��	�,� �pL�g��E��o'�7``Ҿ�6����v1��Xx��TW����c�� ��$�v�b��/S���v,���)��YQI��׍#з�?e��3x�?�9c1f�=qa��rt@�7�\)��éE�/�zS9�p*�Ӏo*����f�!ֱ!�8���0�Y?���/	"=�e��D�fjO�phV|0�-)O-���YSX^X�~�Q��AI�A�ծ
f�1�%�M�