XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����l��;�C�Phh?�u�N���]�|���Ȏ8?`ɣ���!���dtb��{J_�����Bd9Q�����3�〤�ſ��^���=�ņq���-�^*W9���M:����@�]#A70�LY��f�l9��vRdx�V>8��
��7\������MMo�Nb�A��D��<�9Q=
c��"�%��DIa���-��6��ci;	ɲ��.x�l�˚%�@�$S�JT8���-O��Oh>�9�B�=Pޭ>?��!S���|�m�:����`0����Qz�u��F��F������t�B��QN�����٥���N��H�8�s3�w6�]���Z�R����ut>ʕ�D)�W��N�9�
�A(>y�P�p/���q�A@� �c�#W�� ���t�������"��X��m��L`H۽���:�yP��b�@ғW B�v���l����o�8�hCg�Q+�ɦ��gyf:֨v��Z6�/U�FP��}��V����gPՃ�(K�!����q��ȫ�nY����'�����jQuXD���A���a��r�:����c�^���'轇0:���k�/�䎓��<��4>���� ����f��"��s@��9Μ�E��F}w���jD�8��p�{`d�Wk�8+[o*/��^�6���iz}��� ��r^�Jq(Z�7��|Ϥ�Z��\Q|�1�f`��<1�-��`�-E�Տ���mp׸9�ĥ9��XlxVHYEB    41c2     c40MT'����`ql�/���4���s�+{Bw��D�u��,7�*��f��%8�a7��A>$�w�M^!X/��^<l�(Y���|��@iJs���ʻ9{*��-�R������O��mŴ"J�;��%ݴ
��Hɞ�lZ�g���ࣕc�S�f*#� ���vD�	{85�8%,�'�:�PJ=���z��<��ng�ϿHƂF�쮓�	��]�+�����R|��_�|��[�-0����y�GoSJoV�,�Ţp*��z��Gf}`��{�s*�F0�����EM+�x& �*6)�4$s��$�>6�����KhO�<���f<���2��\Px�2��:Ҁ����f�gw�(z�~�o�ւa�-Ⅴf�r}�}�(Y�EUKH!d��;(�O�\B�OL��K���s���0^K��q̹�є��*��f�g���Q��2E��4UkM�]`�h/��[��M�?��!>�V��5Q��n�a�9��п/����c���3�Ї�a.z[��%1�V�I�䭝�s�q��q����f�z5�S@p����>��r���Oמk�̲H���j�fm�ߩ{h	(�ۥ��pA �Ƕߣڧ�;�᧦v���֯�4rdO��K��{��V�C��(\���iB`�ʴ.��/�ym9R������Ҡ�Ij1��B��I�ɬ��ì���s7K}�b���N��ّ���k�<�U�(�ߐT�����0zs��vv=,v���w�������3 ���,e<����nQI�H�qm����e(�\k��`t@v�C<�;�qk���e0�d�Ѩ�E�����	B5��a�����=�Z��n=�=>��z���y�d9L���d�G��}�[���^���)XŰ̂A6��R��31�1QT(�S������K1�V"'<y#�2x;zM���iV<�>�`�g���E3ksM�1M0��r�����J��	��$� ��L��߷$t��e���ygladU�e��uo�.�H�z��~G_��y�j�U?�mK���o΀;���;@�������N���fb�+��7nK��kb�r���4��Ě?{�� K�.M]B�I<D�i��979���q�8��nޔ-� �f�C��>�����(5OJ��%�>Otj��1�"�YL�B�㏏���:���
��\���7_�`?������%�	&�q�OB %�芌C%�To�,��t������Q
 ��7�P��t���o�P7�E����-O��� ���=��`C'U})Z��-b1h�yf�C�{2���.���Τ(cz��6I�p�˼#�+��eSyK�& ��kQ����J��9|xEý�$���t�l����d��O���`%~�D��5���XP�"���+֢aZ�rce]F(&֋H6ǋ�I:�p�����w�3��J�r�2�;-t��3�+
ZJX���(��oo�D�B�� �I��ui
Ef��7����s[O<|:9N�Rl�G���X5fc��y��L8�Wd��ц��O1��N3?(�شv�L�Th�%�*A	llXa=��l2a_?��]vֻ�\��6��ނz+��e]v1^x�#���Th������DS�$�3W�;"Ǒ�*ȫ��1��!��l^eֲ>��G�HU�m��ܲ������M���
5p,hvf��D9�@�=͘8�zp+~D�a�+��ML���^�g17�bZ��@}Xc�	.�_��ծ1 L��:#ژ�}��¶�)�����Fx�̉�lh��4h;�a't�,;��U����ݕ�"���/<#;�m�>?�E���=>��L&�~����6�Ș~yX}?�CC9� $F=/�}֠`��+�|�VɈ|��*�4�W�����)�_�Qc0EG��G�TlB��h6+ˏ*M��!��z1����r��ʴK�ή(v�VS��96>y��FJ�`��7��*��G���Ui��L?q��҃�x����ׄ��^E^R,�@�w3�=X~�DҰ��|�_���������$F�y*�OU���#v�.��H�q�,PLE���Y.��P�o$yӄ��d՛ʹH�>M�m����0�8&�M+
־��V�yy�Cx�TZ�����T.CN}�Rd*��Yޒ��^�.Ύ�D���|�!�"�	+]<��D�@� J���Z��>��l��Q�{���ڢ���'EϽ��6s a�*�;u��.=j��t���zr��|(6u촕%zH��k���Y���C=g��M|�{��x����1b2��o��������t��� �e>�Q�N
*P?�^�t�ͥ��vm���vB�!(��c!+�vi�x1	�e�4+�����ݳ "�T�N9�e �Y<�NLu�c1Ut�<T�ͥUӊ�<.��&�і~&��feXȅ�	M�����J���|�Z�A���r�S��{��0�HyFs���f��>�̝�7��'�<�M?�i��"=:��(�뺄ؐ�c���W`��\N���@* 4H�FF�i��hCH������p�k�}"#/T�d�t;WK��w��{{r<uI��+QE
[��0+����Wo�q?���-����b��
L���H�1B�j��5����8u�@x�J$Ҿ�ZYkJ~*h=�%�r$��ԗ��s�~Kš�����F"��!g����e�{�o�Tmq�˅��b�J�lt�\@rz�ը��w�1�
t��N+�N)��A+�t���aq��ݫ@/���=R�H�``��"����ˍQ�HcY2��b6�,G��A�4����DH@��.��I�AL+'7Rq��>��e���r�J��C���hx��;*����gz��	h��mv��۳�h�Sж�$=O�6���}-�0��"P�5?~���)1�4�m�C�/�6yW�k��9|םt`H����Œa܋����G�ըn���B$1вUl�9HH�-�����x�����c5�G0�ŉ7
t@~���K��/�`�t��*C�#/�2ƛ^`�zO������Z
U��z*�{ ��Sc�:Ľ�K�A�etLZ���ffZ�`�d�