XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��X�D>5ǘ@�)8�8����$Y��(��:̠J8'< �t͊D�/�������P�I<y^gU9h�~�e�����)�i����!U�Mӳ�jN>�3��M�e�/�Š9y��R�~D���ʡ���nyMn��y�j�m�lC��Y{����uT� �xy�:���ꀖR�>Y�-N:|��b���!���l� �Jy�T�nOq�-�mӨ�+�1����j��n(������@g�\xZK.��c*Ϣ6g	[��ZLo��o������C�՜[4���0�H��T�{TQ;��Ɂ҅S���ؒ��������w��f���D_˧���I�W��vΈl�zȾJ�ځ0ܼ�G�Ҏ�!�I�lt �;�d��Q���Q� �i6b+@�Vc!��v��k���=e��`~��7�	saJ̕�C�"Њ٩�oAg�eX!�m����R55ac���K�{E��),�?�q/��4Lv砻�g��t!��`Y"M2��0��p���vLH
�+PS�����pr�Ԑ�f�鍃~���t*R��~�7n�<CN�d�p2����4A����X�)�8yK=u�>M9&f}ۙ$�/�P��;Y?)|�Og~�LC��W'Tk萼�ͦ�;�c�[�Ɠil�x���G���V����?4s�)n�ܮA< w��B�Q��R��m1*�q��@SQ�#[inӱ� ~X#*K��,@8�¥Fbʞ�%� 7!q�.in�Ʀ>6GF���0�����MF�`7g�90�->O�g;��F1�H+�p݊XlxVHYEB     a3a     370�̀����^�kt��mɧР%�����Ԃn_`���sTV�G�w~,�p�\;�M�zQ����,g����Q��/��D��QU�$���Y!{|4�4D1�J��s�ёXBm�=YW�݀ ��<m�k#�t�ɰq;%�ς�ou2�~}漋��r���_?��	&x����ý�Ҽ�l��K��N�B�eB�זUL+��\W�"�����y(�K�ꐺC�$�G�8Bk��`�K7.JHT7��LTHh|�.��\Z�J�M���h�`�h�̧YC 1��uM�?,wX���в�V�`k�
��n�3�:�]�r��)Urq�=S�i� L�!e#ȖQ��-����)����.&����Z�`=�E8P�̑��noȰ�x��a��`=߿l<^u�)V�~}]��]V��=-�χ�yސݹD׌W��-�u���B��* y�D���4���\p!MX�@���ua_.j���촍������kdت��Q�5x�/�嘳�#�S
�G9�z��BY9t!T�,����&�.y9;�W۝c1�~�͹*C[�DC�&�O!Ͽ�k����8y���P���``p�+Ą{K�g;���ٳLDǂ�W۬�]���gm�YV�ƺ�e|��6u����oS��G���.(��PnL���`����8x�%0��O�,�D*��V!*��&y�>�ۜ�D~*�b��(M�Y�N� �}��I��3��@��������ҩ�e��|��B��CG�.@v��4�+I)�<��L�b	N]4G�Σy)S�I���̡�������?�^���B�!m��m��˸�S�RE+�	ӿ��,^o�d�c[iٽ��(s��Q�L�wo���/�%ݽ��>�1�N��}��.�