XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��l 칣cqe(7���l>#�ػ�M��Q2�.\�r��/��p.�=��k��.�~����>��0�@�B "�7����3����GP*�b�i���e�F10�s��r�K ���7�D R�)X_�k�2�1�?���i�[nXW:��Q8錳(��:�������m"�&�d��V���p߻��B����R�DΥ߸	���D$���%P��pI2��T�9�Ce��xW�s�с�C���0s��3ɖ�G�gmf ��)I�h�9	���z��&I�sMeY+pG��֒��{��X���z��a/�=�6��c��3_�EO��0�k�I��A�5��/����0&HBZ�>W/����ER
��D��N�6c�}����&�
�,S�>Z;4R�s�n�q�鞆d�����G=�N�g��g���3�_�#�z7���s��ALG��6b���r3�>��K��}g4��[�>Ͻ_��;�lz��7QF�u��]f���}��iX���n�{�FN��ݴ1|9��YR�%��	�Ƴ�r���]���j�G�Ⓘ�MPÙ�zo�#�T[�f6K�&=ו"���j����@3#�8�n�M7��]���N��U��8��+�ۑ_5`�(ll�J=׽.]+s�n��И�ΒM��a,���z�y�8���?fgzl�k�GU���y-#�Rs栁�k���o�~���c�1�n��B��sf�p�tz.��a���<���[$f�+�z@��XlxVHYEB    3248     9307D�3�~v�ZRgbe@G-p��Uk��H�'-��8���V��8���t�z�(��� �W���P���V��ȼ�%�թL� +�H�0��%�PwBt���^�J��G�;
�u 19l�x�,�j���}c����2����M[w��.�g��X߁u�1����S�v�2D>��4�i�4T�� ��pBKoH����ͦE]��m�]U�/^GGsA�r�~���2;�O��[���,i�9Bu�H�/t� �~D��]z�Ľ� 8%�㮩&������=<��x�I�J5'7-�,k�^�kC�T���~.�P^ߤǂa��b����<L���Sv�Os+�n�L�RS[�p�R��6�
�۹>��L�}Gҧ�b���fF�e�N0��\)~mT������B� [#ۦ�<��a���t�ڽ9_� �VjK�8)qjΖO7����,����2X���T�Z��]�h����yr�@��9mA|��	��qT�6���Z���_��z��"��V�t��@������)� (D�<75�A����|z��L��2�v��թ&�6�ギ�oy�z��0�{׹sG��L��U�v��8��[0+5��E)#� f�ݵ�?�nd1͢Vi�c��s�;nSW	��MbX�6�L�l��g됨�lQ+��:�Y緯{�.
g0h혵-!���6~z�7����.`;�tn������"�Gs���5���T�"�tl��x,'n��y����$(���Z�ʪ*�L��o�NȔ,��_fA�Vc^��|Ve�3��zT*,u�&[���S�(���o��_J+�X�	���&�B�En�y� ������"X�y�O߇��u	a�of6`�~���;��r��e�b����Zi�u̍��ۖD9�S:�xo�/���\_|��.�{ #FP��F�bA�|[y3k���0��X����l/��oo���X�Zs����3Lk�6��6v�iY;��r�9�8po�܍�T2 ��¶��t�� ��.��}�l�?;3��,`!�Ǎ��ש�S9�|U�߯e"l�'��PFcRyd��[�.����v	X>�m@��$��N�d�~E�����xcf��W-�t�s9U�����8���ݔ���[o'ovkY�N `�)SE䢠w0@e��2��Glt�@�� u�����9�-��#�Զi2t_������N���5Gs�lG
(Q�d9�+�\x������	�;ԙ2�ߍ��$�]hbߪ+�%�q�F4��ue��n!C)���2�s�deY����%FvŔPq5���A��&ҏ�c�BC-&֭��e�.C7Ǝ1cXk�I�bĶ�#y�)�<ɰY�»�PIh@r���|�a��*�lrx��.[�r�fR�2�dH�qx�{G!�?�F��߳�lS�3�����-'�[�6���"�.�gFb��`�P�a������3�7��nl`��'E{�Q�� �4}8�[(�B
��jJ�Y�Z�6��l+A��8���n͉u�K[���W�T Oc.���ɇnm��!wŉ�Wow�Ǹ�6���sX��O�$�A�4i�[p5+~rW�XU�2�K�&�ܶ��.��5���@~g�g��cw]�B��G��JnGGs�Y�"���#�k����C�hT�}"p���'H0�9I1S�jO����=��WEIg$�x7�U�sjp1��j��=�u�(u��PF��H2�?F?��������:5�����/�Y�
�1?C��J��wA�]�cɣ����Ma�	�U��ǌ�wd��m���L�՟G�C�iO3X��?Y�����x4��t�?���b?��w�a����Mdn�7�:,���50�,�݉8E�'%��9l,;�Y�Q�ÑKwvי��& A����[K����u��4��B�i�40��, ˒��q�9g��2� wDW����=���w��SIy{����%�����m���t�V��{E婃0
���u��`s�ֺ���G�Pϭ ��NO�p=���؅bX�>�S2,�Q��΢`�?x8�<��sSe�.-���i@��L���P{x�f��&݊.�������s>Z!:^��]X�'����v�!QX���>Om�L�p��7�?���<\��l*:�հ�Rى����S̞G+?E�pb���pf}M���Y����P�����a��œ�r�0����D���^�	*B?ٲ��C�Z��p�1�d##T�iբ�U�#M����L~"w�85�p�-�ʽ�L�~N���?�G����f�R[�2���]�`egK�Y��6�^�0 �n����y�-|I�@�:wޚ{��