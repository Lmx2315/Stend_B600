XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��#=�6�y�
I��%��6P 	"���T�7�����S�C���=�y��,}�d^�g*0/�ر�w���1��̞f��S�F�mN�t���L��
r�9:MM2�Խ8,c�t:n\QD0۸H��Pe
ߋM��������h���3���u�[pbq���(�L�Ӹ+0�1��(���Y�/�'�v�%�ϪάW�w���_��A�Е'7��qr�:ڄ��+H��ʁ:o��<�f�3��qƞ	��L(��v������Ӳ]�(]��;�mUs#f,e�KߥiJ�w�my�MD0ƽ����z~/���/,ٿl��c���=��t7G��p䌕H�����%�UJ_��(F}�Ȍ��q��_Jz�a�ַ�.�YɈ{fu�c!���p C�-`��S7f��I��xmf�;7�JL�F���#��pa�\lJ�l��b��q�A����?IVd��ȇ왠��/`��o���y~� Gu�����BN�f �)R )M`"߾6��\����8�C�g����r"P�[|�u��)���r���mJ�|^�k����1�h�[�;�<R��=��%��T�;�!��^>��'xר!gZ���x�w5xU!�%TY��^.�Pۮ'R�N
s.�^�����b,��*/I���O���۪�Pwm��fu���G"�m�C�ӝ�x��u"���u_��*��@ѶR
���r�R�F7�lf�'i�R�v�S'fpx�b#B#�/'2���K�ػ�|m�� es4nJ�XlxVHYEB    5ff3    1040�?\u�a�r�sʊ���m`b��;D&�8�6Oj�J�v�]z������C�0�'���~� �����9՚�Y���ZU�A$�wn��7�c����נ�u�=]���h�31 ��z%'�
���^�P:�4<���Q�k�R|�̆ű!����J��ƿ-H̢�Kf�i�X�B���yi��6���4mgx�y�68�P��Ǻ�G�i��8��tW�D!�Vēkh��8�"#�& �!����.����Q��Kc�r{�h��߽^]#rʃ��(m-����<�}�%�Yʁλ�!�@��LJ��6��@Oz���ek'�x��85����	�nȠB3�W�f#�ܠ��f�SJH4�����\Q1Կ783BW��hG7�Y �Gl��; �x	s5c�;���,�i��4�
�u�����R3S�ΐ:7^��Z�����Ǒb%���(fq]�YNL`��Z�)�
���2<��9-L\H<y���G�)k��w�+Tn�� ��`w��$�i��͂QC,K@��+����fso��n�^O��m���߯� ��i�]�3|�(k�dxh�k(��Nޝ0]�w~���;+bit�N�0��c���},����르�s}ه99o��'�E�"����_n�V��m���ޢJ��	o4�69<!7D���{)
W�슱�>O'�J��qN�\��1��`cL��%���6	ݭ�/���_$rq�{O�]&L�h�,,�p&n�2v�C��p�Tb�k�'N�v��Æ����J:@cn'8x���i��D�_���b��SB�Pq�������u_pW'
8����ѕ�OE+�/WM�v�M>�e�?T��>�w��ʆ�K�b��.��c���?1T�dF	/ ۾h��Ml#f�`��^����^����y��(�n��p���t�AV0��(iL� l��!�K��$�ԾF'�#��D�Q}�Y�ά>�x�sN��+�S��Ñ�_�r���;)�"�j�[4�bV��Of�&:��`w2�Y��i��&�����a�g���� >ֈ�Ԅ?i���-����,/�v�凄����R��� (��P=����X��zZ]�^С1љ����7ۧ]ȕ���b��-p�V�����.n7	Y���כ���!f�ΐ،��&�߳+���>�Z}&Qc�Du�F�O/ӗ���t��YH����$.�Ӳ+����>i�)A����a��p���?��j��PɊ6����X�㕵U��N-��؁U��9�S3H�mKw9@�j����c�Y�(^����]U��^�	׺Bsm;E`+��w��(ƪ�\�QEF�F]L��K|	��-��6m:���{2�P�J�!�{*Ĺ��/����9�f���~�o\�=��`�6�@�e��O�*v\��g&��r8W�e�����r�X�^�cΗ�4�g
��Q����mɍ53ZV��9٧_=�2��PH'�W ڢ3�S�/�����~��(,W��-���5���JRa��	�Պ�4�ޘ��;�&?��;�w�Yp	N��ֳ78j��֧5s����Ӧo��Y*�LJ��R�NKn����}FФ =z�N8(������h2}��xc0�^�?��8ā[ÌKV�l�����{�j��ڋ��f~Dⱃ{���κ��Hx���v}6q��X՘���
�<��9�-i)Q�؄=+Cd#L%��@���s�.��9Չ*-t�E]ΒjD�=l�bI�2N)��Y3����*�9:���w`ۛ�o�& /�~��Ǥ-0~3���4y��I�4�	j�AXb���w����TU|�G�[:J�g�I!划�����!�y��̸�����	U�S�r�]f��q[��-Kt�먜��f�qb<G���K�����|��פ�R�f1��c$����[N�
��M��:�aM�z��>��,_��ء(D��Ӑ��H�h�[����,{䪧�V:�.g��.���~�?oSK���8c�`�X-��6pAo� ���%I��Q��H��S�PIE��]�>YUJ����j�A�\�,�5�ib���\�P+�:Us����pMo^pRج%b��*�����f��8�YEB����ꥃ���=���G;$׭WU~��P�f�:��;��Tcc�j)�r�u&bt`�J[�Ҭ�B�j��frP�#	�ݱ��`���V�y�Zu��v�E���2ԇ�&%,���#�&6v�\Ii�7w*$�5N���!X�VD�B���ݾ���m�K[�͹7��g)}�SKӥI�/Y��y�G�%\�2�&KQeA^�yj���>A'd�n�E�W��Pf�TR'��.�β B�1��NK�|�ND1���L�f�? r L����Z!x����	��ܳEO�-"�sMm*��ul!�d0�i� �S��!�X����K�����s0	�-R7����� !F	�Я�y�P��?n\�-U��0�F��E�Z}!����\{�F� j��ʮ��ڴ_Nσ}��0�m%{���	c"����Ń��c�7ʆD2kS,[i���e_ck�u{S�nb����Q����47�د�!"��;v��D�9����V�<==B�܅�V���Π͚AmW�ؚ��i-r� �����`�?��4#׆��6���_v�~N���5-FTb�, ��q��� D~+��r˪�Zv�	N��ޜ�l�x�n���E���PV�6t.���+�Q��@c e���� +�l�ء�D08�)�oӫ����wҏ��������#��v��!kE��6����4V�*?�"YF!l���n�&�c�����<���:��/}Iz�]�l�a~�����հ�����Կ+X[6����w�l�I�J~�k}@����#��>�x�x��ᆑ�ZS���&���GI�]i���C��I��Ը����t4��#g(�~�-	���ܦgKZ/� ��e.D �`\!�r2���]��w���^�e%�>��ñ�3SS�SxUU,���(G*�	l`=��Q?j����=��JӚ�B�#���Sr�Y<����.�9E��j
�x�D��l�(5��QL2i��h�uӉ�Q��^Oݱ]ۇE��!��e��ܟ���Lf������:&) aS:�9�W��p�:,�=�N
M��k��i̬�B-��C���T/�����q	�e҅%u�	�<~�}�U���d�{NX�h/<��n���,��|�K���`�(.���_�`n�hcǄ<�n�["�~Xq�x݁���z�*���������y�;��T~�8x�=��OX� -[,M�ӷ�M�$�Q+mq����D��w`G��vϣ��~_9�锶��;��Z)(
����W��v6�d��з3C�*���T�W]"���ٮ�u�u�}]�ܡ��$���=*���_�����og�lM�)��oS��)_//��gGr��ш�wM�g�;�e��������QX���5�8X2��,!	��:����<V��k2(��j_1ES�$��+T|M�P���^���������5gr�h�V�93+�Xvj5�H��5��2R4YOV�`�+�a݀����]���]&8��a�����K(�QVչ:�V�v�����A������G��z�q=ը)�<�C�x��,��^5�Z_ʒ�~A�FD��d.���V�X��4�p����!:�h'���CK �͌���Zy7���"������Ib}=�6�d	���H,2ƣ%��Or�_��}+�_1��bb���15A c˭�GO�ר�gJe�p�>Gh�@�l*�W����!h�����D�X��|FECA�w�بȤV�� }hd�^�U)q既t�l�V�3|nW�m���4�&pb��)�rK�M!����2���<�P���#���ۃY�iH�k�-1K���H�sIϊ�ˮ�:�����@n�b���N����ȣ�֢G��|�V���rAԶG}g���͢�����Jø:<u��O��\�5ظ�z I�ə?����P�.1�D4�h�J�ʟ:�N��6Xޙ�4�踟��x�UA��a�(}�o�rn�e�_"gUC6.gQFVC��;�e