XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���<��祐��x����I#���Hֲ
DM{D�����+B�\(�y��n_��Ē�'�ɜ�mϟ���Kc䶎��H1�S�`��mw�������I�(85i�7��kL�c8�>K�� ]'sߏh$�����p���ur���Ƙ �WJ(��a=z�u9=��`��U";q�8���;�C�R"�R�J�Ag_꓈�ObI� 7�Ѱ����^,G˅^�K؅(6.κ��g���R��#B��f� K��&�S��������r0�;���ހE�1�s�^�8��}�5&2��$A.�J�	y�"���ٗ���	A�5&���6�l�.I������Fӱ�!��8?ݦ�j�~�7�a�| uZ�}�w��Yе����ٰ��b#c�������]�~�Q ja�(��3��(.�L<���cZcTU0�t&�Q�]�%�^��}z���}�Ҭ4�JI����G7�8� ����SY�Rqnԟ�@����P���̬N����C�y�Z�����?9�|Ů�_B&�0@��^��y���t58�cZ�]���]��T�_b�U�t��#_U���/P����N�Q��<�Z�8?O8*��7��̙z�~n;�)
d�`QeD9h("���U�/�(�zU�IDWp{]���֜���)R�fd��_ܻv>H�9l�0����_\9���B0e�^��|����o���_㶭(j�n�P���xHS_2��BS�f.�c�J4���XlxVHYEB    10b5     410� �EU�1r~��%��f���$�~/��#'��4�2	��Q�\���[�%_&��#u)�A�pHe����a��Z���M �d����@�Z>M�}Q���a�?�"�������C]�ň ������[��b1>:���En�M�6�Yw'�Ц�=��uYH���d�(*�X*�Z%%��B�dcϤ&���vג�s�	�N�Q��6~���ph���5��.Z2/�0�W!�y[*:�#��(f�$M�����2Α�����C��݈	�eM喳�c���v5�]��DM����������_��0���1ݷ��k`������"��ޚ�i뤢x�i{���ʥ�oΧ��X�	^���ȹ���8H�}�5N1�����\[,U.)ka��s��,Ӝ��6"�+f�l�|�77�Ɵi������>dl��鵛9��e_�;v� Z����U=��S<��+���C���l	�=^��M�ϐ�5�/��B�,��$���3GY�>�ݔ�f�Ђ9��"�Lr��%�7k��D��g=(f�n?[yl��?���Nm�"����7��(��8V��g�l�UGC��tj����qN���&��&t�_}�+TyBKPG?Ċ*��d2��w����l5
T_��H+v�s5�dk���K�)�D�Ƿ����ϴ�.��ִ�������+#N�keB���<������Ǽ��ʳ�m�Ӕ���1>�\x�ƙkAORW�ֳ�\�X��i9R�d�z����j�4��B��Zf��e�-�mǉ/�eb!%cK'�	1v7��s��tE��؃'��i�Tf7��������,���qZ�'2Q�o�կ��W>_yE�R�����C!3��g�>d-��c9�H�L���%5oF �[������՘�gH��(�����I@#�|�}�,H�Ob��^s��3
c0[�]|�������,�Ä���W������f�؀c&ҁ!�� ��xl�O��c�ؘ=��P�Q�Z�)1RT���h �m b�s��QmLDR�Nx�� ?�