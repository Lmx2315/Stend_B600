XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��i]�g�,���6��ku֎Bf��?jj�6��GZ����/��|>��]�Ym�+ƍ�&q��W����1��e�$��#���xGz���i�$*���tr�w������x7����׭���pl�~Xܽ}��sƜ�w8�)R(u���������
.b�H���x�� ���;��Z �P=�����K!���/�;m�Vq\��鲃�����z�N�Pi::����1�)\S���zFV�P!���[^T�j�0��z3�v���ZTE��ho����Ƈ�/�_��E9v����N�ij�������#3��`)�-K�:X[��]����j����aX�a<&$��+h��?�Oe$���^�B�d��m4����{�򔚥,���}@ƁH����`�gN��O&y=��!��#<��=�?���!�sP�Ȅ�諉������!D6�<�|�>�>�x1
`�H����}1���&��b	��#7�O��屙M�ޢP�O>���������$��Xg|�6'�׺1_ZN�"% ��E���&� �Ǚc��ȫC��ʞ����iJ7��,LJ�0��ݻ�D���U�6p>��I�����t�g�(&Bw]��柋��s�o.w$F�r�7��ɸ�=�Z�H�d����bH������h�� �����)ҿ��-̢R�������:�ux�ϥD �N�o'��}�F�1�N�@L��D�U>RGM~�ƞX�Ϳ�s���Z����(����5j�
��6XlxVHYEB    156c     590��+�&��S�g�V�?�=��l�f%
/Gs�W��+!�;�ZN��BMx����^�N�[���4D�uq��D0SfAN/��M�8F�-�����޶���U ��d::FZ^ޑ�M� ����J��=a�ʷ
l\H]i�_���4�}ño�u�Y-�Μ7ɦȫ 	��'�a��MZ��hw�RU��^�L��Q�~�}�ʰ��zR�0��qJ���� Zns�6�ӫ��[k�W�фQjpI9T����݁Rj����5ef�Vj�J���6}3��F�rI�*J�l�e*���5�!��;<��a�Y�8��u���&(�D�0���[�n%ѐ�*c��E#tQqsOCGB�
)L@-눡�S�{�徘0R�Rڻ��*O۹���'��]l����v�P��>����[BKa{VG��`^>
�A�t�9T�-�R��a��d.�gu��M�}�,�w-=!�v߂<�j3�~��S�"������v2OG�Yn(����r�#���ϝ~��Z/�{)(+�#�O�t�����ߏ�z����sb�Z��M�W�p@I�}�DG��A�[c���Y'���R�E�����;�͌a��Q�#���,�&���l�j���jy�ś��Nv{L&�E�
m��(H�bk>↾�>lM�`�����>��hs�=)]Q��8���im/�g�l[Ag�&�!ۨ��nmMAZ	�]ycj돻��&�[�����4At�U-�?+@�	�ێ8��&�NGX�����4�E����!Z���V{��x9�B���-��uJ�&ӻ���ұ4�t�1���6o�CG{E����8�4	 �b֠���2XW8RpeZ<o}"ܗj:����o�%��Vn ~	pw�7_��D��s�jC
K�@SD\A�z���XV� �wX��C�j���w�Җƽi��EJ���N�+;Ғ(�g�}�a���<K��!��΍�!�����u=|�Ж��k��/>0�; ��ЯO�f���9�qQ�p9�fJ�o��Z{�w�ӜP��Ik�.���D��H�R�ڏ��4|�����L_�3��Ρ���|����#i���>U����p��,�l�+5��s�#z�Ћ���	K�������[��:ݢ���
�����ݫ;ɀAG"J���x-��] p8_�+ K!�
�� D�ش���6��&#��W1�,�h(���^�"C��Gz��J"�êQ_6W�ī�aJ9�~�����1O&�i�|�
)�yՃ�1i�}�&i_�d#'�P�*�gĂu��;h��j�	k	]��].М�(���&�j���Q,���%�f|)xTu�$(��eC�5	�:;r�e�,T4<����i�>n���U�o ��:���>.���8{�����hj}6�i���`�Y��