XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���,F��w	��O�E��p��R��)6NL�n��
� |!T6jDHId�A7U��X�=���~!�/�da����у��̐Ht�ns��pgp�.���1�}�c�*p��RS����X�`�u��1R�ם� �ot�2p��ħ~񼄃q���O��!ܕ��#A _��GW&���t��/�5#��dUk�yڡDJ�DMh��������"<H	W���A!I���9K2�O0��w8�WD%���"�?!�v��>CT`z������a�su���۾mg�[���٣_�O�����º�]������v���KN�
)���}�0&�>�G�/�݃R�� �.�?����E~n��LJ9�n�R�례žQ�����!(L�F8/�icOG���-��e�� ���?2���{�i��π�!��+Bk<u39x��٨��P���S��b�{�P.x�A"��Į
<4�(�c��=b�����C=3x �T�>o�����oe�Ĝ�["�|�8��U�����봆К�qL����a�*}�U�Yo��V������q��=���[�c^DZ-���}�O6���/+=�f[��v��p�2c���0�NNt���hY��<�p�>��	�̙g���T���M��Ҳ˥N�[�ED@�'��w����\)�Q;RXj�
	#kbP?��=&F�����]K��	Jz�޹�He� ��v��R��^h��ngbsu����`֭8�������ri�r(XlxVHYEB     a56     380��%��mG��fx&p�	%��'ޖkR
�ǩ�;\��M䙸����R��Ҝ4Za�m�ߏKǆ��F�T�OE�dq�D�}Lt��[�&�����J ar�{O#�[��nhC�BJ��;*h�e�?��1s�b��Z>�`�B�ϚD�i8m�Y�Z̊�"T�E�9h:r.
��Sw�K��#~�����Ɍ	d�P��8l8De<Y)�Um ��1U�A���*�!������t���Y�y���F���<$@�$PL������6�<YS��u�&j�S���J8��-�md�-9���iT� ۱ft_�vm&��i��W����.,��G���q75LU���WrHEq�Xa���Z�-KC-��#}�Qq<��B'�dpS�	�q����3������o�N�J���y�C�?6k��sՠPMTU]���K0���S0�Cإk�Ӆ��1ks?�-\�TA[w�0ک��"KL�)�,{q"F<�9�K�Bo|T���6t�G���7֘��ڪA���_N�mt袗R �l� �z�Q��]Qk�f� U�R���E50��P�i�i
b�)s,��EU?׉����v�'��������g0؀$��d�����'���ɺtG]&)� �]Ntr�# �}Y��X�pRU��7� ��o�q�x �܂���l�)�C��f��.>(��N�@f���p���D>F�؀�\1�j?/-!:�g|GH���M�M��o5#-�Ku�N��a׌��.�<�Js����1H����D-Ăo���r#��ȣ;f�X�@`�ɶ�郇�
Ё� �ڙ��7p�w����\O�VAOm�{���pv�����������fo�,�N�w\C �g.��*+�ɠ/��e�5