XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��L̂vZa����!{s`d�����YW�΀�����Ң���W}s��6���I�<�Z,+&XnSie�H���I抈���2kkx��lu��X=�?�b{��9\
|hP�!���{팗�܃��#)d<�Ip��dۺ�"~�-�a��������:Cs� J�;��f���#����F�����L���$}���``j?1��3d%ϔ�p4����QE����u{�4G��'/3j{��o_�Τ�0���~� ��g�곦�i��-����.����ɷ9�7������|H��
�g1)
`��O]�8�@4?��ܻ�0I����iX��s��#Q���]v���M3u��cx/e<:L������3�ɀ1�a߽SVc�@��hzLZkU#��h�TG@��0�g�c�Oy������~�� ���/Ƶ#]��]#���VBP�}�*��&t�
�#���K�+�Ƭ�����������3}�ø+���̄<-�V��L����pm�l���x��0k9����!��T���o��UP�3F��������Y[|M��$E��a�jG�����&�R�=� N��!FZ�{�-f5k�f�w������b�|�R���Ni�[6�2j����;���Z�t�FO��]�����Iz���>b�b|�!�BQ�����Ea=�CX7��Id�T�bY�V?�w~��	�s�v�l��zcX��Ə&������+=�Xz]K;yU��? ��XlxVHYEB    3a15     d40���Yq�
�`��5X ����L���lf�b��1r����j�4�N	�A������2���:d��o��fSN��� �du�/VoA�W{G[О2}^M8�LWA��oGu�����́��6��7(�i]�O���=��tw�D����9����GR�/ ]��k��bB�y�Ng��/ �>�v��	k/��գ�ip���L�l��oOZ��S����p���w�C@v޵N��4���}`X�g��iX�ֈU)zЄ,�>�a�H�li��0�
n�5�(��F���q�w
�)}�;2{0R��ruk���D{��`�N��rl�H�E�{�����pxBR�5�ej�+��oX"��K��.T4��e0��1�MY�[p�1&�� 2�<�[�UC^�����;��;��J�B�-¿BV_݈c'�ٕw���͒�Sx|ؼ�$ȍ�	6	�)��|9�O����V�>�r��<F�	�����N��pU��Sk�B������7�4�CY�:D�'�a�,��U
�J��<<�ُ^B�����11pm��m�<�s�*�ۄ0��sJ��t���)4�@��sa�g���(��j�$ް�ԩ�,��]��ȌMѪR�I���յ��Vcu{e瀮2=I?S����j�j��;�
��,�*�0�����.���KU
c�|3����s�;EPS���!.�����4[�*'LTlA�������*y���<�e��x�/ ��5�Bg�HC;�]]^���8�{O9\�<�������r����|�	�q�µ��
������F�&I�����bp>�H ���e�Q��ɘ,TyEn�s�(@� �9 .��*v4��9جro���U4����%�vB�mR)�?U��F�_�,�P='�!�^�`(�Yѩ��VT��n�O���i)�r�j&H�P8-�a<�f&\Ɠڸg�p�~�~7�(�U�B}��lLzwx4^����W����l;JX^uMc&�d�8����e�`�y��]c^�9o[����m��.� v0f��Yw���
���0���n,��1���N=�!��a�t�L��>w��Ru.��[����L�j��`r�0|�蠨]7C�"�C�3���u^�:g�x}�V`�d�ӧȞ�g(�,�zv�M��s�$��ˋ~E[{����/�kS������$'�(q����a@Vm��������?� J�Okm�Ob� �do`�}�V�K�z�U������:�%�et̑�m~S�|YVt*~妔� |��zI�p���]��8�摇�^�[T%����_|^K�m��W�P�j�:��ձ�a��R��	���D��=7�`��NZ��v�sYU�ZN@�=#��S��OK旴$r��X����X/�X��G��BR��Wvuh�6q#,"J�[a��+2��ު r.)��&		�X�t����.�>�W��I��*�(��	z�_���4�8�EY��.5�:��~�L;��( ��a�!!^��qr b�G�}�4Fc5G��M4L�x��б;e�����s#�i+� �V>�M�
70Js���E����\���S�F ��ꪌ���v���LܪP�@��gX�`#dcrv(h�D�8_���R���ʠ���\��1���!,��W��	�#����Jɋ#�co�@u$OV)���4P���|G�V�&��*ly�_��^G���|D��QN��"���|�c5����
,��Xh���ᰲ��rP	��ھ3��
���� _��w�JJZ
| �$Ⱦ��b��]S�f��3#y�7��A� �w�bL���kD�d���%V�1���Ԡfz�lO��e������}R��NPC����?r����]����K�U��.[c��P]��9��i�ȁCʲN1�RȔ�B�q�P=��ֳ��i$A�N�U�:#{��N�Z�Aqi�����A���c��ҽy��:̄v�&��9�~�\�<t��VVjH�ʈ�z�n��a��"*��l ��o]r��1V��s�����uJ���r'�][����>E>�z~�9�G+�l���7�`%U�O��H@�>5��>�Q����)qD�)��i���s�@�A �"�q����K�y���5F�׻�&\FE�$���^cŜ����ğ﹫*�,6RD[	9�Ϸ�����Pk"5�o�>��M\Lv((�$�W����fN9? �Ju�b)�4m^�">�@tˊKHp�l*�o8�gOh|C��)�to����y�rS��X����{�?A#8��r�����'�R�	Q��3���c�?�Nmɡ�p��qVC�W,P�X*��	�c�Q�w�Rl�Ã#@�(b�pu'- ��1�?����Sc���\�:z�v��<0����t�9�+��Q���[0h�ftW}�r:���:�6�ٶ�~������q��@��yG��f%��"�
V��&�6ɜK�(�/�~M$g�E;�Qwy�Q�!6""`~䆰�փ�OV9����b��n"T�6�i�&�����Mu���<߷Z֠�����(-� U����):�~�trv#~�%�mGAG��c�j���O{��6	8&ZJʟ��
�Y���ÿ��Fh�d�09*,պO1�t%(*Ư����_��O"4���$��\=[��# +ϊ�ݵ�=���:s�-�c�S����{�����9��l�Z�K{> ł�d��]�r�˭@&@A ״��]��xgB�=�O[r8������[��V�"#��IR,���a�	�4�$���7��34����H�؊��y��@���������'�b�1k#����釪�����%qY��D�]<B��͖���1-��3,��}=����]��\���~q��^�O�YO���I���Z��k�"I�k��8h�^Έ��D9u�Y�8�`^M��85DbJ�n*m���Rɐ�>	�9��j��\�YͿ�իXpw��`��BM�̈�����a�y�j��ߜ���s�.��N�E�*<�_���k�5qq%��[J޺3J�[ސ4��XX�b8��}R�|�����	 cyV����l�ڵ�Z��r �UKg���H�?�+�YR�'VIK>������J"����^쳕8�D�3N�R�L
�Z5#g'|[�<�5^�M�c\e'w\�^�� y�{�h�Z�h=<����h�HUۡ�\�2?�X��i��e��F��>��J������*�����-�<�YG�6&'8ک�u>M4t�X(%��+�� ��it�|9�fС��Z�Gټ��c�M�%\PA��=M�z)<W�3v�UyZůo�Ċ�Ɋ,o�BL�t/C��!��6��.23�DfVj#=îj�