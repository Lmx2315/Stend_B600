XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����b��l#�fE�I��j �R��P�l}Ga��Րdq�t�'��DM>�)�w^�5�U�6��)��6���+H�	�]�F��`�<��{_�t���WQU�μe��N_���BrY_��D}Gj�����0	��ݒ.gVm�*!���Q�[ϵ}������m�|�����!���i%l�C�At����c��X٫p�Y����R����RWV�E[��!�!�8�Ч:����͹����,X�F(tz6nPn��]Ҁ�x�2�e�	'F^ī��N�/Y{�0��<��Љ�a�O}N=%��3��?�p�}�ז�B���F]�vA�e�m�o)W�(�;�J}��$; ��T��=Z�bYߞ̖�85�L�L�'�(pهK�������{�]Bu���ۜ#h*4d�h����9���6��x,1���	�,%(^�T7=D[��E�<)���%��;Xש�A¿��#�\�Z�
�}�!�܀����������CV��	�-��	�����mZ�7��a
��6fFo����U�>}P�*j�%��j�.8B�$"Qm�!��C7Ǡ�����P<�­�8��:]+[��kY'R���-�K�6�m ��qp�;�W�l��%�6W46�PN:S�Y| ��c/��Y��lX�͢����D�MJ�!��dh�q�[��IJ���bV׃ݣ���N�L���BTܔ[;��Ԙ���D7��^�i兝�n�F�`���3<��9�X�f����2aXlxVHYEB     99f     360�#�~U�b��U ��P�3��0?�k������:� |&�����=[vN�=bDohQ@�HU����2�+hژko�}]bZ+V�+\�"�d�˚���#�����k#� �G0;A�`�昊�	��P2%u�W�_��0إ�l�
����e߶�U�Nnc�MOZT�]�q+�T����4�de.s���0��)�|�`�Z��s#��SC��6F{X���H�)�.|��k�i�%�N:T{f�?3��ϳ@���7�MZ̈�h|��#6Ӄ"�}��QQG̣U�KʧǺ�A݀t���P5�&����]�O|��V���%BC��ǻ��;��,2��X}�4�*t���v[(5{sh�/�p���r2�0e�W	uJ�z�9����9���0��� ��!r7��:nj�[�\T/w*���~����dH�_L�kir��T��e=&���hw��Aĳ��9�*�gD�]"���Ιt9�k� ņ���Q����i�TPBD�ʄ\�oY�%�<
���t ��:�č�3��V�6�b]��+j�J�g��P�vue�/y�5��v��-�[1���.� �T�j�p��	���9�%�g�s9�`i�*|�ĉ�D:֨MR����`�C\��N4ߐ:G�8�<�y�̾�D�]Y��-z(�AprWF��q���Ѫ��d�����\����,F���𳀗�d~-Χ�E�o��&J
$x�bRV����1�f��h�ޕ��ʞ�\~�a�"�u��9.��(�$R}N-�$��ѢI?a�pc?�]{Vq^+K��&1����Jnv��ɪ����z�Mݪ�k�د�~���u�&��}T�?��r���O%t�_�	�j�U��8