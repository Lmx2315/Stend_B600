XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��y	�#����{c��Ѽ�4"�b�@h���<})�%�ކC.kz�,���%j$�m��M��������K�2 �N*ы�I�2�b�l��r�3��0􂥩�9"E��=�sR��e31�|�姮?�SrR�v���� H�R��?�ٌ�s$C-Wm���t��+�`H��[>\��$KZS,;��\t�E߷w��iT#�V��gf,�P��%ǩ��b�V����≧}TmZ�c�yA����ZO'&�D�~��QxQ��m}���U@���P"@3CVh=�K��X���p�J;���Ll���>�@���^H(3�O?>���e�eI�(�.{8��H���«�<����#�8��Ņ�/�������첀��ΫL������1�]L��Af镥�i� ���Y�����)�'�'�ʶ隗�7�M�~��x��\���$����&I�����|�E�̺�G
� o B	��J�M�tt�\
ΔH3T��Iz(�Qn�tU���	�R�4̕����w��i�vt��{�eF��]�xxA|4�C��&�vP���d��;�{ׄ�J˳��>�d���~�j� c��i#Ъ����4�b[W'�J���� t��r�d!G���u��O����nhԫ+ʑ���˕�k�4V��9:ƛz>����:�#P@��TM�Zv���������g�^�`2���q����?����)KD�f��Jy��fd1(� cV�'ɺ?xD%�XlxVHYEB    1044     4a0'���=����y�Ҡ0�;��
� �R6��c����ZJәh��ْL�I��*��u�(�'L'T�Ous�o2�#�Y|S�jc��J���>�X����)�����I��ѹ�ğ��GP��m�:�}I��FpK����1=
�Ou��{�����i��Ç�-��xOJ���%ȑ��D߻Kq�LJ��\��6�j~���1^9I�2����L�ˌ����k�>:��X�m�]O�x��5�1Hw�K�p�H�04�����jQu�~q�][+��#����Za
�O}�(��3�Y�!�X,��)��g8�a#j�B�$R��<Z�Mآ��dzj���Ȼ
��|㮣���]�T`���,L�	��k�<�jWB/]<�Y�%����}�#'"��(d���B�xgW����l�4Nt��ч�)x?ϟWm�G��ݪ��J�=�^��8�O�.��b�1$tJC�PHW�����ш�>ك|8�iܸ��jP�`���#�L�*ݏ�}7�.��{�No\V�Q������H6�zC`x��O�r{�&4I=��"Fl+
�VL�%Ų�'O���Z;��[@�7-��@��D����Ul�N��jƘ#��-˩��A��/] ���	r�4�íe0
�`Sǈ�``3$M���nv�]S+����:��4�E�40ʭ=��?j<'�c����u��V�L�Z�,6��:!#��v;�Lb�I�y^q����֏=Pa*��8��t`)Jg��R)�����3D,毫Y�q����k��&ѓG�׫�Yڻ4��N�ؗ� �2����@0P�2�(@���>��ªQH2LY��>�C߷[cj2��;��R�������(��������&yȃ�-��PW���qzW2�H�We���SJ�bpt��Э�l9�%��)Y��Ǚ�*~A��I���l���O�{��E��1q�#H�e\!�����I)+k���{¬ClƧ�Uq�ZX3���憎v�2���-�V^���D��d��?5�8�0���w�ܦ���tɡ$*�H�Oo�3��:_�*�4 k�h�f�N������9� ���~s��`Uܶ��ۢR��u;m��K_� �`���$�]���� ����|�d�L˭�d�ohmM��|����.g��v�7?f2���y�Q�+u�#�/3