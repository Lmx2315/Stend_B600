XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��7Ԭ�,��=�ֻ��S�'�M�ԑYJ�r"�^v���O�Oz)�pE��o�8
�b�����u�Y|�Ы ����9�ww�&+Gcl��������n���v�������㨉�+���N}�9Q�*pI�	��WLo�$*�Pep)8 ߯Lf���$KE�̡�;���#s[E�|��}ui;�>�n�#�Ⅳ�v5�e�+mM��o=��
��u�vVQْ=�E+�:t_����4�|]�A�c�V�#Hk���ʙ�/)�!�R`ҁ�J_}GHTR&�����+���?�K�m|��'E��(J��+R�v��m��+�>����?������	����D���EbMV�����6Ŀãx$��J�%B�2vS����b3���(͜�<8�XA'n߄���pG�|Yj��,��ac�K����6s-m�G.���ɞ�]H�ܚ_�e	�-&/9����f�da"M}�]�����i�p��J����_ktwz��⪐"� �d����q��~�����	��pH��/���Q&��2dwҖ���v8��?j�mAjmQ3|�%a�#$�_����S���9�G$h�����4A��=DD)�M��W��ME>�i���R�Ļ}��t�"|x��O������J}@��H؉��ߒ~� !ȫ]�7��Y��g}�����;���{/½�y�� y��pk"��؅��~�&ms�v��6^x��poaYS{�a�pA��[��|�0�V�O!�Y������!�V�j�XlxVHYEB     ab5     420[D���c׎2��js��.��/gO#WFr9�I_)u�i��@���2Έ�C�с��%{�~(�al`���������H��Eq8H��	���~��[m��:��قA|
wX��[ꃁ+ڰ@-��E�C�Z��1z.�$N���\8i�<}y֡=�"���F�H;;��yR����ޡ gޗb��;�(B�b���r��I�
S��d ���FZ�du¦��x΅jbP!�Sx�{x�;�x����qxy��9�y5�>YO32��qh�~@L4�uH��Q�n�-����323Ԑv=��8$��H�b�T`T>�`X$"{0.H�@�P>�	[�l�$rn��_��L8钢�[V�f�z�
����f�h^c��g-���Z��A)�s�ﺈ�"�tcd��4a+fD�v-�{N<�"�.C�/���;���ɲ������X:�$��1�*l�Z?���y�SÖ�B��YO��������?7�X��o�q��m>�vš����?��W�N�ʰV��;�����I-�7�iS�ѧ�X)����y`�T�'�qr�Tq4�9���R���w��"����؁~�,e}ڂ�)�7�;S�?��״���o�ڹ�qv���"yB0/�-	,_���$i�>�BB�>��������x��K�[��e��PY.�yZ�M�N�֕��y\�uG"֔���>45m�"�_ABjO;7���o�$6�o*y|���5*�����@�~;����1���{�Dª����Ϋ��`�wC�%= �̌mp@��De}���%ȍ
-7����<ãa�4QPž�����.V��>�������磊�j|��|	x���*.\8�'$���?�'#(�[[It����0zTo��r#�fis'�]~�K
!̭�����2Sӟ�C���I�y�Q�k�f6,�˓�/MKh�����J�p5�f�V��k���[�4����8t��Y�5�E�"��3�����Î�+#����z�Ζd�P5=�!	͡k@�
�cZ:���3���+f8�F�Ά�0
"p��F��