XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������u��W9l�#��f]w�j��l-���M�?�1��P{U�����f�߿[�Ͷ�>{��O��ŭ�ТY�<1 &b5�A� ��d�1���j�v��l���
X�R�wH�������jh���-?�w�Q"��_��[���db�0�h��!?]Ȕm�aѕ��:�@j��I��ث�"�[��\0�uQ��]�g9J�5yp�n��,�t��E�:喞��V���=��:�#<�AЪ}�����-�{�V=fn���Ƙ	�S7�q�\�M6�QZ�8�{�_�ȟ��a7K�Z�X��Wڽx��'�����v���4y�EtX�� ���8���[,r���c�N�5o���5�6�*���5f����y��v�0@�o(����p�T-,��-�X}"R��6�y�����>ڞ	��-ngﯞGxM������gW��q����AVc�o�s:��lƟ,�1���v����h �T���|H���ѿA!1�
������\�=*�F$F��N��Hz�"0b+�d
*��Zʃnqgh�ט�w���A��k9'��?�(�d��B�%�f�#a�,Y��8�
�8ɥ��u(�L�AT���$�����A���+�oTt�%E���u�D�I��g�Y���rA.O�|�,k.�#"~�?���ț<XT_ >焤�D�Z6O w7�0_;��3�������f�K�4x��]E�I��N*��]�)��b0L%J�&�F���8�ՌXlxVHYEB    1cf8     790L[�j�zฺ�������]���a�Y<��۰����S}!���9��U��!f*FPR�"��tiU�v���@v�v�q����2������4���p���a�|bGȒO��Դ0��������
;��H=p��������|���i��ZdRw������=��k�Ϯe���C�(��ۼp�EҀ�UuԌ�j)`Ge��&ޖ4�T8�UQ�۵�ץs�y��bl���6Xk���JeH2T���j}t'2��Z�Db`��a� ť.�d��+���L5>�<�c�}D���~�����,=���7c�o��X�_��0��ْ��I�@B&�V_ˍ��d���n,مT/n�S�QЗ�F�q���m�����WߟEGyS�vACS,��ڪ����r�=ݢm�Wů�&t�����8��	���ˣ'�v����R��O̥�ۋ0�|�E>ߴ�]TmZX����<�/�?EA/�E�CH|�DE�тvP��������w�Sz�J&@�����(�s��u
S󡨧\���h�`�\�5�/������M6 ����Rz�AȔ磬]��c!��x*�$E&y�:4Y���|b?����ja��ïe�=�1p���[��iU�4��$こޥ�B�6���:��ƒ��G~T�v�*������Cv�@�1��tTR^7<y�1�7s�n�"�%tq��h�z�n�6Tq����Ր�\�,�.�رBQj�<�3Rm��=�������9��#_^|�"�QR��=�)�N�_��#0�����&�� ǥ�~���1��/��ψ����MZ���҆�?�?�Q��h�����IO�j�nY���c�,A'���].�2=�P�%x��l��َ�]s%�+��'�AjK�S㎣{~�0	z�Ѷ>��KR;�*�e��6J	y$_�=*�S5���S[rSY~��.�dđy�%�3��˔鿘w�DCG�����IÃ���c6��С+�rE��*P��2��j�Hp�P���^l<ûG�O%5�y��>�z�痍'#���;��~?��3^B��j-iS��k�}�%��M��r�E� 2 Ӎ��jS�c����M�l�	୚,�e���7�)NLh��<��{��}Km��D0O
��XP4ԘK͵�=}ӋX[�Fx8��j<W���~#��}h"�Y��P�&�S�m���A�-��iɒg,������a|v��S{� 1�9�(��ap�m���;�BYdjL׾�8��d{�����.�ں�3�~bJMrV~ׯ�)5�*^L|�v��W�ݪu^O����L��kT�F*� �-J��+���3��d�.d||�P�|��[�^b���6�Ϋ�����{��J����d����"�Q8�|��*�F�$
��7)��~���(�U�<�I{0�� � ��ٴ�/d�98��AL�۟�w��C��j�� �}7�`�P;}`��(�QAjzb���	�M�h`�y��b,�nX6U��\Bn����W>� ˧�^�[�K�г<Yg��o4��Ka�X3A��vZA�W7��7E>��Q��j�2�fE���6����Y�~!�6`+�'�Dt]��mm���uof��_��G��/�f݀9g6�'h�.�r34M�?���>+����cF�t��b�X涜$D��o�gO'y �9�wV]��8��ʻ����̌AV��t�rWvzq��W�Ҝ�c_��հsp�K�쉴7�8N��{uƯ��[��Uv��l����������Lm��=�	����|������\L�>& ��o�DF��[�0&[nIM���g��E�m��<L@�P���F�]S�3y���:_+�ɢS����ͯ.�9��Cx���e^�|�J&���A|���T�g�sW����a)��̵�0�88�%V�