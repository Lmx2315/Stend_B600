XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��JZK��@��0�f�2�c��R�L��;:�H2��XzA�ߟn��O]Fm�g�\횅�� ��` U����!��R�X�nw�)����Z�;�R�����߁&%��b`����0��=����_V�!<W+���p��a�h��C���i�o˦G��&�����/D�_��Q�u�s��J�c����[	g���s�n f�l/K/�wZu8��4.����?j��Х���'(8`�W���}M�i�����s+��7Dr+�;]5Q��K�ْI�[�)��u�@ۓ3ɇ���=>�����~��k�\���W��S��1R�u$wYe���^�Z�sNxd�,�I۸�:W�*j������Q��/m��6��h�?���<i��KmS/�y4�)FͱY��L!�dd�Rk�Ҫ��*;~����Ϛo-���k��o�ZPg�0�)Cs��������*���TN��#y��W��M���&O�S~j=��W�̇��L�b{R[��M�k�ط{}@,	l�	b��!|��׋6_f���ttM��5A6�K�M��;���ߏ������0ԁ0;u������{�C�E��:yX%(=yS�I��TN~�X�+C2���,��9���:D������>6�ضϰ>�Vg�o�W����%3�͕�9�X��$ML��/�9�ZFA<BPY����LV�{@ U#L3ո܃eoS
�tt+q�ów,v���D���Y��+�m-����XlxVHYEB    26ec     8e0��,��At5���"c�nAG
������y��x�L/����Ӯ <z�I6��9���~�E�� �bzG�'�&S.P����%d�b�ժS�	)|�"��Y5axR9�!BKg�3�]b�A?:�*e̿Ōuǝd�+���`��TN��pBc�;�� �b����K �5wK�������f���)�PC]QLH�*CNz>���\J=)�Ҧ׸�Z��jB4�њ�D>���}N���X��P�A�-���[��B F�  ��'���� ^�
13SB����0�rk�ۏu������|����J�EA��>�9�k,��6U�81�������1�8�H��'j�a��"]N\�I� v� I^���/�C� �W�y�>8��t��c?q��h�z�R���m����_`��������L,��LƦ�6�5�8�4֦�q�F��&��0�\�⃢*�I��eo[��V����.�ו�����"n��G7l�." Kn��{½�w�O�Ȼ=?�2�����z�OW'
!�������,�}
�β)�h��͓�,�'���.h�7S��g]-+,8�m �0]8�yNj$�7����*5N��@3Ɠ��N�=�(ؙe-LJǴ��]�z���-�ݽ"���к��It����Ьw��gU���m��"F�p5&^�h%�#���Z��;R+M�7'�&9QN�C"I���ݿ�W���Z��q%*��Ep�:�V��9�
$���{���ݓ�m�Z
Sޅ�.P�d_H�or��J���z4��I��1�,��^:�I I<Ȇ{�/�V�	�gw:!�s��:��r����E&2�
�J	��k�)����g���`�m@a
�N�XRj��I��4��T��W^�%�����c�/�e��������Y
tǑ9<MSV%K  �Hk��sD��[8�Й!�DuXk��f���5t�V4I:���g�;!pƐ5^���&��Ũ�Bg��tA�0�Qr�c-��"`{V�L��P��"B|ؔ�v:Fxx�V�\���6�@�Ls�Ƞ�(����Ե�Y�A��H�S��=%z-+%�O���C 1�B�5��K��s���F��@�r�ig䪈�>M�8����KW�\<k�L�+`a!je�8~!n�=V9�;^���]ƴ�I��qW^�Ѫ`�*��������G}���cЀN�}���X
	wvn�7i��c���K��Z(�J�w�4Z��������>ZZ����Ŋ���-k����v���@y'_8�=���ZH�ʲzrĆn�h���Źq�k���f���➜'�ġ�{i���𬿑���FqT�Q�cx��I*O�Δ�ȫ�M�,&�"r�`hyƐ�]��uO��('{\�h�]�d�&�%��z�"�������~�-� 췼�n��⃧k~���1��{�G�����O��i�y��`OH�M�Xǳ���ߵ�	���?%��)\a�_�A�2ە���ķ�����y�ڡ.O5�TL��˥X�p!w�5�=�:T*q����#Q3{���2��C�DW��q�Q�Re��	��v0�l k�4����������Fv���c.�$�h��7��􊯟� ��'CT��Ϝ��hf?�%��C% G�&���?ܠ��{���=U�ЋX$��hA��Hg��k0q���S�sa�`��Q������.k��%���y�����`n�.`���5���e<���5���<�Xy��/5�_�[/�3xR����?n"�]�!/ ����k����|���c]��3���P�$ B��>�����C�ˇ��b>�?��RDH�#y���̎�3��Hׄ�'����x�!Z���ª|iN�_��&fsN�!�g�����x\��~)�#ǂ�:�`��-;��5##��O���K��{O�^]�C�pp�= �PPa�a�#7-�¦"���Jl&�7&�3�s�Qm*9��a����q�3��-��ᯘ���ZSP��4��nY�hI�8&�ht,܁�h�z|ff7lPf�m���>)�z7Xp�E.P��%'[J��d]gC��}Y�>&�BW��r�J�<��Ԉ�Í���
F95@�V,�X�M�;sU�H��D-;�CJ���O���g�@��	�>(�tw��c���.cq�F;�D�uH�O�?��"[���-���ꍞ��%�A�;��V��R#�KɁ�ؘ�3�X��ό