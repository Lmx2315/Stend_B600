XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��V�V�H��"S��&�S�6��5 Q���;����'7� �e����I�6��{��1\�1n8#�qk���L�V�63�nNUĔ6�������P f%:�ؤT�Z���)S	�Q��T@^�-�l��LJ��=o��\�4�Ӟ�=-���&l?*��ά���p���F�w���ӵ��B���?������֦�����C�2|x3�qt���v����©+%�������L�0<#��:�'<��"�S�D�/���O��	@�Y�aC�?:�K��^|�K[a��rĴ^EhN���:�ԞqS��_�5� �w��@{W� �9+'��N���l�с��e���D"q��	�����!� <�W�]5�ϐ��i�lNO=4�D�e?�_�����;��@̃
5�zЃ���RY��L*Lڲɹ�~�s+9�֋�%� ��݀�P_��- U�� a��2����k&�-�t�;�:A�~�f��ئ��?�OX;�q��D��
8����':��_-HR�������!�Z��F����X^�	�u)ͪ`�e�,�d�&��=7"�u���q��ȧLX6�^ۋ7㣞2·��$_2w͸u��.1�����37]we���F�~��H�#B�fύ� �y;��ј]����_�]�F��?+�<��|��m9Ϻ2?T�gi������	7xr�T����)��j֭ļ~����X*y�V��/s�FcJ�~��;��7s�	Kl�i����_c���XlxVHYEB    7a0a     c10|�-���<)0R�,ȓ#�Ԧ���Z�Ő��sˊ��K��]S{��v����t!ɯ��<?���/5�%F�8L�HL�#c4��s�N��+)���R���ǙG�H�P�J���j���w���<	Cz�5������1�Yy�:bt�*���@�]��ix��4�HI}�)�5���|��{_S�kKz�r]U�.�:�f��`��NR�3�������#���z��-O�tU��T�@�c��:�-(�#C{��ZUK�0�𰌁*�<�*a#�c�����/�V3��L4��������Bì\��W'oP���k*�9��X�t	,�ݿ�
�z6��|?tz{"lI˛l�����b�����z����(�/�@�ѢMU���FU�M1H�V���q��&���͔?�E癤b�*K�L�;x��g�<b`7��?�wcr^��5FBVn�Ac[aƩ�0KK�$*;8� ��*�"��<S���.�o:�Y{nx�ͱȐ�f{n2�zF��F�ޜC'M�2[�}��SѫF�����6�|�fὉv$�O�g|����y���c��!���Y1pAmk�T�/Q�
gi[�J3#bk�:���Ӌڕ?-H�<o��*�, x��]���.��qT^��Οw4�e�ͳ:�B�O8ylV�n�����y��P#K#5�1%���w	Pۥ�Sc��J��Y�M.6���'�ddN,��ܢ��<T@�Zc��B��b	(�WP��V�̛���;M5k�_#�O~�v�~�mI<���{c�&�0l���Y�{x�{~wa�y�
�;A���+5e��HH/��
�������&�)��$NQ�U@�}?��7㒧�z�rRsn�8sL-Y��)}��N��`��e�]A�����>�1��]F�ZXm�*�ꚮ�L4�h�A)�e�hÂ ����lTZؖ�,Tbq\��@.k/��Vp 4}����T�N�Sx�_��"-V�|���\�+2y 7����2��]�����w�֐PQg�	��B}x����U�;���Y{2����Ưv�Jy��@i���fAA�E�3^9j�b!پ�<�^���<�PL�v��/�zǃ��z��_;#W���A�jc BmY�uİ����B��~�0囡�f5HX9ܶ�h��A���-7��qXs��6��7���>�h�+(s>�ޟ�[i�)c$J�0����jL����k�{�^�U��^-S�?��_ST2$�
�zP�wW	�vO`��:?�1Ǧ���LIJ9�E��WNPK�@1T� �-1A���L��3�����im�Z�{>S�y܃���-�ߩ>�9��7�ٌ�'�0s�o*�ޔST��Tl�6zs�;�Ϩ�S�e�|3�� 8c�"E������}]�}ËP�
�������;׆g�!j��a���|��@��8�]fg#Z)]�d����,�m��p��U�C�.�1' j�����~��,|�cg=X�TU*��$\��{Ce����e���	�
)����3~���A%O^��z�Up	�iݏ.Ȼ�|%�Z���j[_������w5��s�.��h�S�~���R�Dյ���Ó?��F���ýҀͪvI�|�j�lV�+a)p�,'���>�J넚����Qȳ�n#7��?!����Zۤ�(1��i��YA~jč�j�iַ��V8��i5o?HD�ز��&k=�3=��ɉ`�m�Q�]��yi}Nv)Z&��%��nX~�MP�e�p�^�l��
�g���aH,ʠ�d�����00N�� c]½K�<G��}�׮|
��b{���?���j}�lX�`t%��{`ſ�A��9��I��A*2?�K@v��<w{�h֧?�LT�q�[�o��9�?B�����:���E��( #��]OʑP����c¢�SN���K�/|>خ��L 4s6�����y������&(��!��ٍ��h_��j�:�T�S��e��y��+-Zߒ�[�j 9N=,�pw�N!��|�p��U1��&!�z �(R��B-m=�I	��y2ĵ�X������@!Y��"<	��$H����Ɣ�OԞ��^m��7�� �%"Qp�~ʜd�:�55h٭�����:J������2).����R�̄2=����,=8q��i"���cy����]���/�e'�vH"?xY!�����?�D�,}b���a���^Tg�mt��u�0A�>�mr�ɶ*��6&���]c$o�o=�GT\���x�T~Ý<r��������K�Y�����D�vg�Ń�����ZT����U]�~�C��:+�YM1�V�eA(�L�׺�� |��3��A��oN�{���+-��9�D���*_,~+X�\�|@���#<~�09T�f��tΤJ}��!�ɂK��9coe���7�W[��gy�y���/T@��5�+h"�?�Ji-*��5���;ȖC7.6��L"*v^��-��u�$��-�t��� ��-s��c}YN!�����k�0���r��ܝ��M ��p�\7Z�9%�&�	$^�R7I����-	���u~t���X�aD��
ً3������Y��4	ȟ�t�u��6X<���A��Jq���,B��#ʁ ������6�=+y* ���X�Wf	T[���R�}�!� �(�h�g5�Bҟ��À'����͗�zD�όx�L�A�I�K���$�w'F���7�[5�i�խ�IB ���wS�*Ո«م6��9B��֫~$QKg�c��QS-:��hh+��l
�Lt�5�����ʛ<��� �L�<!�p+��og��Bu�CJu�p%���{Q#\�����H��I����ն��AvR�g՝N�6}����.��m�"]p�,:�j�v�Bn\Q�K�%�k�[��j>���yѵ��mbgN�0|�d����7mj�=����`҄2<'���h��՜%����w+;3cE
�E�e���<d�\��uwu.���q�%��B�Xv#
t��������5y�r�wi�>�]�