XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���=��(�s��%C[�������a/&��L�'PRy�/�u�ŏ�͚���2�j�xG����������b��"!��1i ��n�����G��P&7,J3H�׋�ԇ58��Hݡ�\Ǯ���|�%��s��"�ͣ�k ��̔͋�Cn�$4��Ҝ��_>)J��K&���8�rѦ�����6�P �$+��h��2�0�̳��$��0|Ɔ�(YV�/��Fk���M�ȑ��xS ���
n*m��5_}����-�s.q%>����<�#MOě"fd�C�3���D��30��R�����U�`&��I)�BA�l���Nu������+���R�W���U����,��M�)�8�ӂ]�~���g��FMO����[�HClr: �0(�J���ݔ3�0�>K�, +Ȱ�ZB���>�5��S"n���țp�|ح�%Z���7�JƁ��xNF���d�8P�jލ�!���|��|7���$[ڤ�j6�PZ����<���}�0%	7��+=��ϸ��3p8��� ������Н�)=l��@4�3�P��\T��_t��J�dpK2Z���]S���w��p�y;�z2sIՈq��M������%����8ga��)K}`Ec�dg|�7�?��T��HD��'ݷ������͐&�ДuPj�f��N�F�$�NE
��9K��S+�xto���m=�(
O���- �M���q�ĕ�gK�?Q`+���"�c�djm�e~�9�+XlxVHYEB     82a     300{�����O���wE��a�%[~ۻ�
���qw]��<��sex5�@��L�~� 3�C�JR��ST�ȴ���y� ����c0��NG�E��﬐,6¾vw�&��'.�(����Q�� �ѓ�!6��eU�K"ė�3n �)��]|j�9kG鉤'+�SA��n��D�� ���sV�}Y���A!2gӆ|SE5q�����q���<K�(ya�C�̭ޝ�#s����x�*0�\��J� �� <��65I���( 2���|ʾt(�[�;0%�,X.����:x���k��M���SY��Ŗi/[�2Z���}��<���f�Z�q��1���K�^f�
V��/;Wc��f>��!��� B�[�S�ކ.��(�pT�6n�.puɢ[ E�l�	��S��s����)��e��M�p���#9I�')r��> ���[�cv�~<W�&�s
���Q����>�㞯K���}��:��0�+v)��#�
�oӂ�P�1���(B.̵��t�V��0g�V��I�=f��e�0�:^a�ugI.�篽�}�L��)��>e/����^>����8��Q�m��fr���� d`�q,�Y/�B�UϘv�m�>���b��]j!��Z훴���	P������MKXh��L�Mi��5��걟�1���Q|FaI�ǅ�B1���&�H�d�:a�
m�X�9��/mcpyZ?�j-��󤧧 �ֶ�n�u���h����H���|u���c�E