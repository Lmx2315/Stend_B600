XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��=g6��C%[��^���j��/�K�l�ʬ�����8GC,��'��[�:�{qؽ���b���jW��^	ɏ��n��(Ϥ�x4=m�-�+�5�j���u�FH/�Ɣ�%e�}��1.L|7q���vT�Od��YQ-c�]�G��)_�^۳�X��%jMw���Bm���@c�#bnf"n�xAR(���L���q�Tw���f,MI3̓ްp��=�?q���D��;5o"de�F�
�2nõ]�A���9ij����/o#"O���=��fU��W�+llI͛Ӛ ��Ğe~�`�`��l������.~�R=iz�T��t�o���~��]���[�go�Z�)�!���@�*�@���ٱ�l��IԀ�
&~�w3�PIHf���s_e+R�ø����0���H*�'��L��蹊vw���9f�}�.O�s	5Tw��,1�A�Q0��@t*?tGW��x;a�*
�������7+��1�P���r����7�H�ch��@ D+�$�O��\iq�P�'^z�E�ۗ�Gc#V³�Q]��so�TGܢ�>�<R@�OK���$��?�k��OhD�b�I8�&M�6��$\������I�v�3�0���`�� �F�F�g��a��K0u.o	����S���65�8�T|˭��u�k*ޥ��Ӷ����u#j������B��;�A�]w����f�1�Qx��4��ϰW�_f�,�Y0��]��=��~XlxVHYEB    6df0     b60�<N�؈�gR������<�`ٶ�پk�m���ŏř1����u"}2�ܪfSo����9S'i��a'����7�y4m�g=ʍKB�|'��Yy��s8d�,�[�Sc�D�ԨvLn���P�~;��Sv\�u_�s���>5PI�0�*Ɛ��n��m��i&R>N*�.��� R��Nڛ7&B04H�t�Q�"����)�%uŵ��}}5�b���"ϛVE:��zs�m�{,�l� �&�q�׼�6���G	!�|} f�����q��d�z��/����=kN1{��ƣ�deM���au�h0�����]��L53�,,��7��uhc埔^��j��R�9e��A@fgl�ÍO<]�ޞ���X�^Ť�s�Ok��i������~k��b�U�,O���O99�\��µ"΅S^r`v��K)����`Y#�01H ��?�3]'�&��v}?�2�{gҾ��pQ*1��ڝ���u )���Rk�>G��s
)�(�_ni������� ���K���ed#������n���m}�e�r�|����5���я0���r���N.<�����z_xB�x3e
�k[��}��Sx�c���z�;��t�x��VR�#{�����g#��m]soɯ�kFB�%����m9�g�&T�G��åZ��|_��Qí��e���^#*ůB��Y-�e�@p���ѫiM~�<<�MHh2��	jh����sM⍏��Y����o��{x����L-��
�A�D�Θ8K�w�u�%�/%a�i$ru��>j�~�����5���9�&�0���ޠo(� &��'x@�����eIcX�ʼ��ΰ}AS��L�A���zV�gѼd 7^:_msrF��H�?�4���=|�f�B���dDN��t]?��G�Z��H�4�&��wqyƄ����ѵ��x��8EI����0��qK���[�;�� fv �e��MspW"����WeH�[8�s�h#��d<�����ģ�.`�O$�ý��>��j��� �w�v�=۔��E��5ʚoas3C.�IH*�(�v�ΒT
Z5�c�����.X�O�M����I_���ş5Q.>�)�Th���h�
�22A~�
ۘ�Z@�̌)��.������"o�Ь�}���E㽨e����&ns�];)Fw�n����Ð�SC��K'��P.�5S�,�|�[H#%�^pE����<��x�4��*�>$;U��/��Q~�@����g�UG��WeTl��>E��=��;�EJ�s���,��%J�'�$�J�����л���	�b6eMX�҆]ޓo-1=����X�4n1M��t%��:+��r�z[a
g���Չ��7��+�{�&uRl���h��hA��6x1woӥ?�>ty�Q3-��s��2݅ӟ髐��/����lZZ3�i-q����(�gGb���n5�uX�r�Xǂ�;��v[Qj��:�I����Iu����t�\X� 2窱Mg��p XU7��(K�/���h0�W@��y��Sw\�Ʈ�Y^B��S	'�6��V���$�vϼ
K�$���o�F�Ж��J^��VMl�����u_`��9g)�!mT �p.�n���z��=�¾�#Q�k<���NY{N�yOgs�$a�C�
>�)����i|���0���)��Fm6��� Ш&v���[�Oľ|��l=��T��j�(e�ۨ�q��m�Xe?���?�e
�@3E[CQ7��A�UQ��$E�,�1�RPFS�RH[2\��S����7Pz^��,���m�=A��9��D����Dc'ʴ�*�^�z�s���t2�c���@�fqa�>i�q��`6b,���_�_��ͮOX�N�Bbj�[���w�����=�������pe�nq�+ѩk��H�F�8�m㩉�MJ��)�[,l���#�?��N|N~�f76Fp)�#��YWP�0y�!f����%k2ѽH]���%v��-n>���nP�,/����9m�e�V<	�4����F�]�β�Fy�*�lQ����NM
->�)�ڏ{�'�*W�R:�M�ǐr:�`�����ɗ*��������iC
�>�z&��$7��y�ώe`if�+9h��{��_i��yd� �48����9?3eNa��J+BHXFP��;H�]����C����]��>Iހض��]�Th=�}ݥݟ�EB�c��K����*I����t�,m�Cc����M�M 	��&2d4�
�oJ��Z�����7�_kKM���aAǰ��\�����V�=M����X��|������e}��
"ca�ՙ�O��쑲��RF�"q�"'R��V?C���ŋCe���%�\�ݯ��/[=~_^��"�p��V���K�dd�������w|�pCT:ݢ"�m����O8�b���,u/��A�N�ۮ3v^o|��^��v��&��+!��n��S�F��U���f���` ��U@[�b=]�5��JD�+� &OR_(Ɲ��W=A�+�{>�j�5��m��P��;<,���dfbF=�(���uX�v1�gS��O!���8b�_Mi�o��S��D�sxjMz
��[�H4\3�E#��#G� ۟�䁪�x���ӧW�M+���}��1I��$m ����Ţq�G�Tc8j<I�D�M�#0�}۲t�T�ȭŴU=�${u	~��p��PG<bg�<��@PP*7��"Z��e8Ʈ����l�͟�b�ÐJDH��M�k!�;#~l�9,Y���G����>�FW��X��~s)/d1v�ɦ��$h��U@U@���զ"{M]C}�B:f ���hn
T\��"�q��#��歷a_8�qa�ks�Y�nk3�U@=:�p�6c~�`�ݴ�p�y��[���Ai��0�[�R��+�Z�C