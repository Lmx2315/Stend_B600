XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����s#|1�4��"�Y�2�q�F��a+^��5����{���1��=^ޅ�5�t��/����̵HX�d0Q�\�vJf��r�Ι�j��+vT��D��3�k^'�*��V���/��߄�oY��"%�5�� B�J�����?�vߒe�f��|U�w]��͑�fI����˓��{K�G��;�7��s��q@g�?c�$�c�"�h�rg�7�k�'7�#�oű�
]W=�y�I6,APV���1�ge��b�}{O���n6�[�"j�	��+I��Zz��`��({oIA�(�
6�r2H%����ʙ��'�GΊS���A@ȁC�6�K�}c�����������Q���� �a���z�}�tp�~7�EW1B���@�6��x��%�y�BZ�YM��zIv�#������5��^ĭQod��w-����乆�U��ӢSc�i�Im������&w��!!�X�2��M����]�"���aL�z�Z�HH]E�G�ӕ���)���C��b�{�G�<Ôf�2�5{�JkBj��`��a}����IH%����GCC��*r7)$�M��M�q�\����~���!�h�'2�K^���b��h��|��o�=w��&�Q�g�&�����N)���C�+J�>�g�r���&i�m?�M��E)_���܋�w}�޾M��5��](���&ש�&�"�k�*�w1�v ����,�����^�UU�?��±O�(ݫ���C�/�]��rXlxVHYEB     9cb     230�ݪ��+,�C�Y��	kI
������"X���>}�y�r{/�� ��E�wǤޓ�z������L��gC0"8��r�'����>�� �������^��;bBcD��@�g�- �6�q^�z���L��b6��fF�x;+&w�q��_ٛ��2��v���	�F� ������ʷ?Hb��CR����`��xHMM��ɪ�K�U��TE|8���E�Y���¥I%wnX��a�A��?�H0ȽMOM.v
)q֣\mR��leR�=�pyD4��ě1Zj���;kK<+�5�|�Y�5�lM!è�PP�Ƽ�U�Y��u��ذC�"�I_D�T�U��Grk��h�j�
����]����#�4̢C�y@3�ns�%ݔ��./��3]�"�ʽ+�M:J�K��	Asa��{��/?�@�~�^��P���6i���<"j�t?�7�3��%LQ��V��<��4�g�wF�+��,���!�4�4?�Z�T��V~�P�������v�v�>�Y�Gfr�ى;�����H}��Y&�.Bb�O��