XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ߤ�`2�_1�dN�����1��#1x�>D
gh��5���FH3�{lMLrF�N�W"�b���=e�$^\l�f��;��JT~/\�-R�g�u�]�4��k�����Z�a��G����ʙ���l"�fX������ K&`y���ȏ�Z�v��$�iq�d��>�P�.&��ԚI��k��'����w2�{ �ս7�_�Ј%>Ϋ�-��������h�>�ފ/+��s���e����8��ݲ��Ûm SbQ�ɽ�V=E��5{��1!���ek��@a�6L�Ȭa}��Oa���C��g�V���h��@YTu���C���:�� ���u��66�b�FS}�l�����|N~�r���/�O�0�o̵��f��@��j�7vX��9�t�?��Q��'���i�_��w� Bs.��/d��!,e�@P&ٜ�k뗨-�A)�c�@~$R�
�w:<g���JȲzQj�����7nbn��<�cj!R�؜�s�?_��� P�'�8�P~H��Z�am��'$hn�p���<�����@�`�]�Hp�.*��q�p3���	M���a� :Z���[B���swk{��E>o�U��%BVH��iĿ�y�0�dV������ףE޲�O#�<�(u q�����w�ǝU�$���x�*�g�N�2[�E]�A�u#O�Z��V�en���5ĺ*[BK�*A�A�����D�GdNw[λ��N�p���i�F�k�7ʂ�������/�tS�����&XlxVHYEB    1d53     7b0xa����lɶ��#�IS�8����������5���q��*�A�ٓ��������6%�Z�v�������n�nrL�<�ɱ䋘�Zw� �����$���e]<5Yn~�J�>*����;ZSGF~V�����NAL��5�au� 7�)߬�aۍ��{^;���������6I罣���XJgY��ϝ�w�c��=B-)D��^����#u�M��ΟȵG>���}���]q>K�+�u?^���?���x_G9�*�$nB����D&z��~ęg��硘�]A��i/��*8D�X_ݒ����X�@�L�l�)��yq�c$�cBf,����
����o��x���(�̙�l�3��	;U[D��I�l3�0A���������0u��&qyڹHm��tu��7pQ��bJ8�[���ك-ѳA#S�Ʊ�ݻ�/�6��㲲G�h�bϿ�fhNϒʲB<�����B�Đt���t����՞|�ol��޿#"\�>��yL�\��b���14�.���8;�)*s\x�uvF�(uz����q٘�!n�&4,]j�S/�r=b,�r�>�SO��ݲ�m��oj&�I�c2���PU]�
Y���V馮��M�V�z~nc�7=o3�"���ug�	��q-0!�c�8�5r�i�%����W�]�Ch��t���)C]	g0��WR��kpы���(S�%�e�i�9�T5h���C�x�ƫ�M�VR��40����)�2���P��F��M��88����@����-��5^�β@Ikg���:���9z���$A)n��f��8���8�M��� �[.)Y ��� FɃme�nq$[FP�ҁ<��eOE���� ��S^���}���r���Y3����\�����/:��A8:m�@�hO��%��ٔ��x��r&6����@c��jd��V��aV�!�v"�\���]dJ�/JĒ�K �ϗ�<
Wėt�&� ǁ��k�εg�8ſ��k�[�_�U
 n�<q��~e���l9c�|XaW�}kӑmKP���s���L�_P}I�*���$k�(۽��ڏG�d4�/Y��Q�*���U`���؝g��S�z��<R�mw��� m[��\F�K���˲�Wy^k�j������YAEn��W�?o�F"���O�Ep��`9�߀�ol��A��
E��9��cB�T���!�v_�Q�6��ԑ}�rk��ҫ[⾍!n]��LiԴ��Π�n��|�
�KStlF�lq�����"�U:��C2���O|�B�b3�Z]��XMף�`�XG�c"�����@�|�foA��+<ٖ�'p�j	��gj�kG_p>����!FC�1�����,K��m��_�[A��i�_l���/!�efis����ŋ^��#N2)QV];��&~���=��O�m\{�#$G�3Gl�C��q�����3U%J��=i$ݽă��қ�g�x]*lzB�:%y�U&�C�1������ޟc�����䖯T˝�Ԯ�l��r��5i��M�a0�T����&���yɄ�)�2�]�����+��%������1�����)MU$A�-�wU>����W�7jl���d��<���[�e��tZ�t��Q��O��!�	�����4�0��\z�6�D%δ��V�GT�!*q#j��} C'#5އ�XT���/aGU�0¬��7��z��TY�>����s�G@�"��妊B��D2S�%��y
!��:�	s{�j�w��v'�$4�˫B*�[O�(2ƥw�\q�6n�:H��-��)���b�՞���4/�~��'������{����>WA�	�S2ώ�T#���4x���g��)��.�8�Qг�`��ѩ�.	,3�Gq^;��7����|��q�S�?�%٭z�)vQW[�