XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��r�j�b�L2d``- �IY<��B�V��܌!b�;��t�ţ�^^bq�����/Ex��|�VB���~Q�LK�B�q�<Fw@h�W�&����UA�c����2�Q�r�����}}��\b�y�r*��]Uh	�t��+����������Yu� 1�{��N�#�����s���0d��Ah�Y��%��yyI���8\W�],�0r��ˠ=s�=Ѧ���>j����e^c����h8G���,����cy���q�$W��,���@��]6xֶ�N�%��<L!`�{�Xjˆ��Cꃐ3�{���������Ԓ m	��G��ogHv}�d:ov�q�2�h��U5�9�=��nc��z��1�*,{�%W� 0�ԥ��Y��1eN`aX�x�g�(8�Hr֞G��'�֊	��L�>�j���@Cؗ2�\Qd���f�w#4Wp��ӆ��A|%��̱� �C�S�X�Ǐ�có`���̭�PP��1I�h��_���n����UZO�L*4���Vl�SP���^��,ʵ��@�n?C����<�CG�g[�6�I(�Z�bl�T6������5I����^���m��i�N�QT�UP�9�{�#��8���x���Ҫ��kN�$��A�;>�͉���ͧ�CI���զw�Њ�U/��yn��L}��=��wG�藁1���0��=�d��b�ΊH��6x�s�a�+����P�}q��L�XG�IHyޙ��˪��In�ggd�^�^��%��/�XlxVHYEB    5ff4    1040�,�d+-��T1�s�ng�������I�Ez�+ܯ'�'s���}G1r'�i�X����Þ)7��"_�MWdB�I?��6TF�p�� i��t����F��2R(�߆|#���r}Mm�-h��p���ך�ڃM����a	,���qf:G�-�\L_[�7��������������N����_j� �����lf��d��N������#�a&���}-x�R�ջf�D2�\D	�X{|M���Y�V4���_#���N��D����e>�7���1�3�r�����%h�2�Vy�W���������UG�2�&d�fXK�P9M�p�ʹ�H���M�el���m�*I�M�Dbe�v�V:�u��P���Դp��zQ���#cA�}�V�L�O;���`-��!MK�I��ϻ�8̶9�K*��I���@[��@ �?@D[0��O�T�(q�c�ݦ+�!{��i!�/�����Ճ��)�+��B+�S-�`���I�̦�pWwF^��Pv���NN�{�#��4�<r�x��Ѓ�3����YsK&�pI��l��61���NM��G7����H�#���We��K��c���K[��۽������Uq1fԨ�}���uM��d� �����5�B�x�P���MOWCz���4�� |B�L�:���Q.]���=h�s�pԃI�ИJ�JW��p�K�p.�c5�C�	�3�ǩs�1tc�$=�ۨ�
^��:h�8fr�� ��nx)O'�]8��e���7�u@3�C�<�ಁ(��yM�:]F�x�@�b��j���!+�̔�kicF�6�^�	�fi�&���Dc0'%r:ՇQ:[#�?�U�A���0%�v����Rw݂|w�(��2ѾG~�0V�Z�&rl(-�����vA_�L����	��H����V������H͋��<����VPv��`u=�����r\�<~&��O�"�O���f�h`4 ��"hi��
u��p���~_݂�a���ۭ�~V�%����@����穌�tЖ��4@�Fl2�$��^�$�R憓^<�T7�״{Kn�(,���)�!���;�)��X<�}���v�37s5�$�1@�QP.�+Lz����O�+�c�@н)+fo��vf�GՋlg��>𖜋�<��1'��z��� �+p�IG�$w��+�by����)�y?���s>�G�^�g�썬��!������o�����/ݞܡ8	G||�҉���V\NpnxR��M4�vZ>ply���ěznX��;ݱ86��^5 �D��Ơ�H���l�}L3>��J�%�v�Y���:�Ozy���d�$�5��<����7�J�F�pR)Df��8����h���\g�!$/x��h���q�mE��0���D;�hqP�.����U�g���P���!T�"�t.-��ӵ
���[�&�>�Tù�׫�U�����.:U+��$�$��  E�E�J��YYo�׸��Q�*5�0���\Ӓ}�=�&��G"-dt��]Ӟ�mfʺ�x���:�]�h����	��h k�� 	Sɓ//`:�=�	�KL~�";7+cS�w�.�/�]��JfJ�6��)���z�u�2�ϟ�DB�R�GySG[{�`�#�2�g{�7�7,Zӝ�4���`�)Q��D��-P����M& af��8+I/..��0�b��T�fy'Wi:�ޕ��II'So�0���@Sؒ��-g�>�P��<!#$Q�����˪�Q/����W�\VۃZ_�>�~�)	�{�zNS�'�����P��Sax���b�� c	k���1� ���9�|�lc�0־��ψ�_������Ѽ#&�O�5��$��GC�,F֌��<��`��'HK��y%`Z��/�h5�<~���4������7��#����6�dP��T+5��±�����.�ⱛ@ȟ�����Э]�X�~�5]}�Ej2}N�ץ�����ǎ����p�)��:�qA����i�q��J�v)��&������qh^`�����J0�a0r��%�'o{܎�����1|�-�d���1���h���v�2�.���.�zTkl�W���G;A������L4d���#[�_d��va$��
�bX�o@�>8���(J��k�juF��X���|o|�߬����%�������9E�B�#{Ց�a�@�-~�3h�( ��b� ��Iq� q��p���;)RBG�(��p��1�$M�u����}���.NV�c�i��$����-��E��I�A�^�9�|��&�����p��˴���� _�;7�k�>�e�x���E�DOaW�ÊN���?��x��Y; �/`Dg���$��r��n%~�HG�:��SK���d�7Q�>_g@B�+\���x�z����7��tߤ�!���Qy�1�.�Iw���25g8Y|���C��z�hh}h��g�ΌO��eU��	��p��D
��Yi�gp�3+M��4pﳐjY^����SXɖ��$��3�o����h}�-Sc�ydK�����u����k%Ҥ~�4`��W�M |����k�耷��Q𧷹�̡����9!�k�;@���7o}}/�ܱ��l��;2���],���h�d7JC�����X�j��V��`/�%��n�i@�8O&6��Y�H�5]�v(`0}�k���z���l��43J���Ruh�{R 6y� �%��\�{1��@cg� k������l���ٜ"�+��b�/�$·cX�o�w%�y(����P���wK0�'�e_- 9D2p'��z��a_�wPۙ?Ŝ�k��`�@��؋ f���Y�P�'�Ed0����UurF6!K1ײf���hǭ0$׫�w�wZ�i^�~�����Ő�x1N���l���]�/���H�_��4L�VuVv+���Q�5�(c73��m�#S�Q$��ϝv��[�6e��{���]d�'�����7�ƽV���@_��B!C+��'�ԽQ� �4b�TI�����?��Xާ�a��%�5+`�%Zr���|<r JíEd����.6h$`��C��2L����iR�!�����"Z]@��;��:���&̿�}dG��V%��Z��v��~'2�f�����~~�g�S)�&Z������t@%=� 'ɂw/80�w=�9�I$��뙐�f?h��8iS�<M.q@$0k��c��XS�F~Lc���	y$+]�G��-��p��]VNH�`r�COF�'�)o<�{{R�"��Ǆ�y�iwV�l�O�߄E�*};�Q]��ޤO@�	�-�~>��l�ُ�7��}��!��w��o��;_���ߜ�T��͋ϼ�_�L�p]Dky,�zy?h��Z��=%�����Z.D�<7"x�.(L�q9��e�r�kr\/:���4���M��5���Ȣa���P4-n���?3_��b�`�^�ȴF)W��%+���o�����˛N�H���*O�5�b("��=�0�@G�(�Te�WS���Xb��|@7~|0o����#��H+�k;?��	�(w���t�Frm��dل��i��5�rZŘ����D��J�u4ؾG�T�'U1��b��mj1��ys�����a^p���5��7Y'���]����{����ub@əd
s�ѕ��`Âa��k,�D����O�s:Qj��w�_/��-����5nԺ 0 X��i?4��|�:ư���"�A�X�n���8P����\�\o/��ߚ�>�O�������Ρ�xXg�Q`{�Z���N�A��\���K�>ױ��6�W���^��/tY[t��Q���8P������m,vy#�BfI��� )V.,����6P�I�թ� �vߙ�$i��tj0����Q���(�~��},�6���*��U����"���Sa�o���_w[�ԙ,+�GBw�Ķ[Vk8��RQ�I�����"�(x���@���4Z�mY�bs��c��>D�F��YUc>���z��ri�Ij���*��_.���z��n��̶B[S�����;mJ[Y�����X�f��:�C7H>�!N+
�T�.����vC�oBTz!F����$b�9q�0�V)d���