				   			 									   //-----------------------------------------------------------------------------
//
// Title       : WINDOW_TRNG
// Design      : DSP_180210
// Author      : User
// Company     : d
//
//-----------------------------------------------------------------------------
//
// File        : WINDOW_TRNG.v
// Generated   : Fri Apr 30 22:40:34 2010
// From        : interface description file
// By          : Itf2Vhdl ver. 1.21
//
//-----------------------------------------------------------------------------
//
// Description : 
//
//-----------------------------------------------------------------------------
`timescale 1 ns / 1 ps

//{{ Section below this comment is automatically maintained
//   and may be overwritten
//{module {WINDOW_TRNG}}
module win_sin ( in12,clk ,addr ,out12,rst,rsto,start,starto );

output [11:0] out12 ;
wire [11:0] out12 ;

input clk;
wire clk; 

input rst;
wire rst;

input start;
wire start;

output rsto;
wire rsto;

output starto;
wire starto;

input [11:0] in12 ;
wire [11:0] in12 ;

input [11:0] addr ;
wire [11:0] addr ; 

	
reg [11:0] a;
reg [27:0] S;
reg [15:0] Q;  	

reg [27:0] sr;
reg [6:0] addr_l;

reg r1,r2,r3;
reg st1,st2,st3;


assign out12=sr[27:16];	

assign rsto=r2;
assign starto=st2;

always @(posedge clk)
	begin
		
		r1<=rst;
		r2<=r1;
		r3<=r2;
		st1<=start;	
		st2<=st1;
		st3<=st2;
		a<=in12;	
	   addr_l<=addr[6:0];   
		
	end	
	
always @(posedge clk)
	sr<=S;
	

always @(in12)  
begin 	
		
S<=a*Q;	 

case (addr_l) 
			0  : Q <= 16'd0;
			1  : Q <= 16'd1621;
			2  : Q <= 16'd3241;
			3  : Q <= 16'd4859;
			4  : Q <= 16'd6474;
			5  : Q <= 16'd8085;
			6  : Q <= 16'd9691;
			7  : Q <= 16'd11290;
			8  : Q <= 16'd12880;
			9  : Q <= 16'd14470;
			10 : Q <= 16'd16050;
			11 : Q <= 16'd17610;
			12 : Q <= 16'd19170;
			13 : Q <= 16'd20710;
			14 : Q <= 16'd22250;
			15 : Q <= 16'd23760;
			16 : Q <= 16'd25270;
			17 : Q <= 16'd26750;
			18 : Q <= 16'd28230;
			19 : Q <= 16'd29680;
			20 : Q <= 16'd31120;
			21 : Q <= 16'd32530;
			22 : Q <= 16'd33930;
			23 : Q <= 16'd35310;
			24 : Q <= 16'd36660;
			25 : Q <= 16'd37990;
			26 : Q <= 16'd39300;
			27 : Q <= 16'd40590;
			28 : Q <= 16'd41850;
			29 : Q <= 16'd43080;
			30 : Q <= 16'd44290;
			31 : Q <= 16'd45470;
			32 : Q <= 16'd46630;
			33 : Q <= 16'd47750;
			34 : Q <= 16'd48850;
			35 : Q <= 16'd49910;
			36 : Q <= 16'd50950;
			37 : Q <= 16'd51950;
			38 : Q <= 16'd52920;
			39 : Q <= 16'd53860;
			40 : Q <= 16'd54770;
			41 : Q <= 16'd55640;
			42 : Q <= 16'd56480;
			43 : Q <= 16'd57290;
			44 : Q <= 16'd58060;
			45 : Q <= 16'd58790;
			46 : Q <= 16'd59490;
			47 : Q <= 16'd60150; 
			48 : Q <= 16'd60780;
			49 : Q <= 16'd61370;
			50 : Q <= 16'd61920;
			51 : Q <= 16'd62430;
			52 : Q <= 16'd62900;
			53 : Q <= 16'd63340;
			54 : Q <= 16'd63730;
			55 : Q <= 16'd64090;
			56 : Q <= 16'd64410;
			57 : Q <= 16'd64690;
			58 : Q <= 16'd64930;
			59 : Q <= 16'd65130;
			60 : Q <= 16'd65290;
			61 : Q <= 16'd65410;
			62 : Q <= 16'd65490;
			63 : Q <= 16'd65530;
			64 : Q <= 16'd65530;
			65 : Q <= 16'd65490;
			66 : Q <= 16'd65410;
			67 : Q <= 16'd65290;
			68 : Q <= 16'd65130;
			69 : Q <= 16'd64930;
			70 : Q <= 16'd64690;
			71 : Q <= 16'd64410;
			72 : Q <= 16'd64090;
			73 : Q <= 16'd63730;
			74 : Q <= 16'd63340;
			75 : Q <= 16'd62900;
			76 : Q <= 16'd62430;
			77 : Q <= 16'd61920;
			78 : Q <= 16'd61370;
			79 : Q <= 16'd60780;
			80 : Q <= 16'd60150;
			81 : Q <= 16'd59490;
			82 : Q <= 16'd58790;
			83 : Q <= 16'd58060;
			84 : Q <= 16'd57290;
			85 : Q <= 16'd56480;
			86 : Q <= 16'd55640;
			87 : Q <= 16'd54770;
			88 : Q <= 16'd53860;
			89 : Q <= 16'd52920;
			90 : Q <= 16'd51950;
			91 : Q <= 16'd50950;
			92 : Q <= 16'd49910;
			93 : Q <= 16'd48850;
			94 : Q <= 16'd47750;
			95 : Q <= 16'd46630;
			96 : Q <= 16'd45470;
			97 : Q <= 16'd44290;
			98 : Q <= 16'd43080;
			99 : Q <= 16'd41850;
			100 : Q <=16'd40590;
			101 : Q <=16'd39300;
			102: Q <= 16'd37990;
			103: Q <= 16'd36660;
			104: Q <= 16'd35310;
			105: Q <= 16'd33930;
			106: Q <= 16'd32530;
			107: Q <= 16'd31120;
			108: Q <= 16'd29680;
			109: Q <= 16'd28230;
			110: Q <= 16'd26750;
			111: Q <= 16'd25270;
			112: Q <= 16'd23760;
			113: Q <= 16'd22250;
			114: Q <= 16'd20710;
			115: Q <= 16'd19170;
			116: Q <= 16'd17610;
			117: Q <= 16'd16050;
			118: Q <= 16'd14470;
			119: Q <= 16'd12880;
			120: Q <= 16'd11290;
			121: Q <= 16'd9691;
			122: Q <= 16'd8085;
			123: Q <= 16'd6474;
			124: Q <= 16'd4859;
			125: Q <= 16'd3241;
			126: Q <= 16'd1621;
			127: Q <= 16'd0;
			default : Q <= 16'd0;
		endcase      
   end             
                   
endmodule          
                 