XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��gtA�o4�I�%�3h?-8.��V��F$��GuN
��~B�.��T-�� �x~L��*�g����c^�;/{Mx"s+�	��>�K��lb��v��cҦU���i�-y\hyy��׌�!��IA�(^h��zH*�U������Rdz�z=9�!e�8��a�xB��E�ؙ,ƭ���ȡ9̠����SqB���Umڔ%��	2tx�3TǄ`"��m���%������/&���H���|\�M����'E���a�~{��ܤ�*I�i�s�ͶN�Z�KKvP���+Bg�x1���P���?Ҁ�h�ϕ��y�Ξ@��p�v�<u6��'
Mɀʐ�L�S�oQ�[H�g�p_��p=��5���w�tVD8X��g��Pz�"�(X)�%%��������c�fT��� ��u�糏 9~�=��ъ�� ƚ�3��͌��R>hGl�t'��*��{˫^�����b�$=�s���2Ӝ�qY��8�Eި��,�|����{��D�(�^lu���l�.�h5=�u�%!�"1o��ү.�����צ�R��'�:Uc��	\w��h.��F>B�qC=�ג�V��gb��ax�b
����g7���f:}.����5��L�=�_���_
�r/~�9�rX��N��Z/ْpR{�L�]�n�=Ő�8��,T��rY���������:KIT��X}ŷ*�w=�H��$'� ���~�|��d:E�0hNv%EB�e$G�4BVXlxVHYEB     b8b     3b0�f�)���`CZ	+6��A��S��CO�@��� y!�e���<�T��}�~�4�L���T1-�JSL���H�+!��W��1~=C��4L�?��]��+���
���IR�B��	^N��%�i[m&t�^�֗���M(܂�����N��T0�������Ԕ��T43�Bl6�9`Wڇ@�6��=/��w����s��3F�t"]4E/��6�IM����.�ַ}���§'���ۓD�t>�q��/q�j�1k��K6g��}����È(D8���H���mF�~�{�dVB�(����ٵ��=�K��a-jv�{M���+I��}%�p$�`ԗ�\ ��1���dH�8_��>G����b1R~Xʹ V��8��#L�fH�V�i
o���٬��(-!]3���e?�E����0p��ʠ��Z�}
���Z=����I�4�ړ��;3XM��k�J�hՔ����`e#��,^HG�̀d��t�9t�:{�~CJ �Ce��9�K�ˑ^=������o����D�"�/d,#򩏖Q�N}��	���_�^�֤|�c×�
��X�N��42��V��ӣ�ׇ�ɶ��¦7����C���/X^ �[λ�@p�ȴ���wk��z�x�#�$���K/��i����6���)nx�Ac���َE���i�KA�I
�7�.Q{�㙘Ƴ�v�k}a��|<WW���= �F���v�K}N}�؅=2"��+�GטgT
 D\W%�ݍ��q��ir^uy��ܤ�#�[�h�Pi<�le���W������4XQ��:��%�u����W]Ш�����E�g๎5��X�	8f8�7kͽ\ԨC!}^дl
�7���M����^S��Z�R�KZM&�]����[�����)��QG�ӕ�t�:���D