XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������E���=����{�4�<�㓮����(1���(�M1�h|f����7�b��<�H�^���A+�?�?~Y����C�g����ȸ�6����c�}�E�Oc��Ҷ�k�ZL�%t�����ڠ�vU�&�el����l�e����Kh�$���{l�5��C"УJV�Ђ��O��
|���|�3h������Ӱ�f�R��Ս�C^��٤q�N\_"��3*~b@UCg��̌�=n��9p��V ����fw2��A8��0 %Q���ۖ��
��g\ݐ�G�|,��O�����d�UDS��LlE��(���B[?�E��_�rx��s�"�x��<�q� p��"���'���*�񦬔�щ�|K�K��(�vn�[�X�)��oˊyQ����ۿ���k��^:�gQ�b�Q۟ʽ�=����S��.;�e�Y�p�';9�W�3�a���j�y6���� �.�Y��)�����J*��V�����2,F��t�q1'P���%�([elڳX�Sc��#فZ�ɴ=M|~s	j34R�HSo.A�3К�+$u��$a�X�u��ƅ�Ή���)����/	n�a}�_����7�0)����@�����UT�%�<�Ų�����k�*3���
H6��os� 3�ͣ@�d��v*a�+F�`�ͯ�i��`߈����CS��K��������]��G~DI��X���?�G���#�o�/��4�T~�f�a8�C�J�<_�A"�AXlxVHYEB    156c     5903��	Ż+w~��Yh>]��Z�9��8W�b��JF~j�l��9}E(_s�hEfs��^�H8X��F��uh�����n>�T�nV֣Sb���UL�{�3=�����+6ʘ�/!��+$�L��4���Ɖ�j)�#�>�m��q�{(��NZ��Jja��̒��
d;�ȓZ���8�2S /t#"bX���3�R>��r�2�9�aRv)��*-��/]�3��e	b���#��-��A� %a3�L®��t�'w��/]UE"P6��x�쉽������e/IY+g,�Ϛ��(�d<s��N�������QX��Â	`�8�OY��q��*\��d��v����KWD�4/�prta�ݡ'K1I��G�"#01D+�2��#�նO?l����ʚ��df���|��XVu%8���sHj��t�<�������MY��Q�FJ�٧�'UٔA��k/�kJ���25d�E�%�C��Ű�2|Zz�����<���2�����/�TZ-�@��bL1��>�y�"���]��U}!���`�=@a!0d���Zʴ���������}A"T,B$8jlI����P�  Όv�U5a�����{0/��в��8U�Ѕ#����G�2��)�m#��*I����!Tt��cr�z��R��� ˺@@<�:O�:7��`9B��n s�|r:m�k��)K��B��CR�@��N��-�i�Cl%ބ�@�"�y|�9��AiG�H{�Ȗ_��?#��^�F�Zj# �� �R��O�=<��_�4��ɽz��|7%�c�n�_��"�{y@n������(�/Z�8egW����<�s:���R�� v�2��
u$76v/��D2�mx�+�)<�%)�g��_�.�����k�d�i�$��u��-øyCʹ����ޮ��A��y�Z���^�N�W19� ��!5wXg	$�4�5�r�S||�݆D����'�E�G��o�"������w�6���9s��L~��;�����f��N�k�2vut�O�'�(��L���u�v(*�) \ ����I=QA��<��$;g�+%�ڢU���.z�L�,@0M��irJb� t)�<I�@���&4\��R)���P���c6����5=�Bt��C�&��T�U�w$M�F�]X&�Y�:���hD5b2u�"&�;��@�V���נ�߯�A��=B��;m���S��L����=؎�d�i��g��x(�_`�b���'�:�g�(��Y��+��
27������l�I��D
w4=;Sn�V�k&v~|@�b�������+��$���-D��t�C���*ԧ�f�������l�r	��<>�L��kE�}��G�2�x��zZ=