XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����e)"��y�)L��B�`T�P�:��z���.�d���. ��LoHz�0��nGL�/���0ԚI�\B��2��Rl����WM��Q�o?<�t�p�,� �:���!�Q�$H�{#���
.�b�%��s�4#7.\ߨ����O�#���f���G��=4��=�҄�&���PyZڟ`��
v)ˠ��A�o��>�gn[�#)Q
�uUgP�X F�de�P�c�#ҬN��,�06�'�Y�%3�#ϣ=U���޺������FǬ�ӊ��r��u��p�/��.i����E�
��hPG�;"������iƭ͇��J�A!X�bn�������٩�t2Iv�՝_R��f2��E^�����N����=�!r���eM?�k�<���z{d�^(�6�ЦX�:Q�W�L��/���Ub6���W�5��s����Ia�Y���s�g0��kF�y�H�P�ʑ%Mo>m�x����{���yN;�
e���4�����=��VSdM�Lm��h�筘�c�Y���C�w��!�w�l+��y��B:�����v��/j'�/ҏ4�[.�Xd�st�����[Ud��ЯIRzS���qʙ��(.�>F}��Y�, R�������eH�F�.���k/o0���)�Q�0�e^����}U��3���D��s7�&mV3�k�m��!93۱�q�y	��[�{�G���RZĦJ&M�E�Cԃ�]!�/
P�K�OZ��.V�{/��c�Oa�G�H%�8XlxVHYEB    3c90     900tZ'����c��BH�޼���lpU3R\�K/&���6�ם�%x%5�n=�;- �����(ք����x�<:����x5o_�&��p��?PJ�i	�U���3�2�ٲnJ�d���[�/��'�.�%�(�?n�_'T�,J^�%b�YYa����h���z�������������#(n������*-p�dK_����7p&�]���^���^(���id����� � 5ó���"�5�x�K4�D��%�+f�\�|���
��SsǮ̵�� �9�<��/���Z�~-��g�.MG�V�)��Hz��2Ц��D�)��n�xp,yyjO�o��is
��8�� =�����-������� ��O"�1Z`�Bb�_eԀ𠗟R��j_^�q5���Y�A|�Q1��
p��]È/��ҹ�v���'��5s��ݭ �uCl�F��"H�qAD�r��fu��+&�����\�sFu�+�.�"�g�_��أ4�[���Q;#,2Xoj
�ױ�O?n��.��t�C�kƩXY��ß��	egW�s&� �[�j){Z�O�d��3��wȰ����!EϨ���nN�qp�R��'[�|�%�4��D�Eq�V��n�iD·��y�nz����
�3E7�+Si�t����K�?Q�*���G��,4�ғ��V�p6��v��0�5�W���K!�=�AC��F��%�ty&~R�e��S|�ft��e��4e���?���a�ʾ2-�9�u������3Y�
�
�i+����U�qv	�u��ȚȬҿR�o퀄b����r5��� �3��ҝqȢ�آ�vߌ9�^�R=�x>Ĩ��!�1��q�u�]r������p��ۊ���A{^'��`2�@��X�=S��G)v[f�$�R51�����1)k�9��"�,�y�Åc:���H���p佷�c։��kb�=&ws�Ρ�f�K�"����+v�ֈfv,��[CBC��ك8ug6�����aG�[Z��ص2�=�����j#�u�/�b~#�7�%`��Ql8#�(@�Xum�e���h&�6�^g����ݽη���c����_|�|�\�b���u�-EJ�������98�k�#-~4>(hoz�q6�m�����d�u�7�/��8�g������ �45�Lꎋ8�WD��C"�)�j`y���Q�W�*�^��<tJi�D ���ܺ��&�����@�OѠ��Ԋ�����FM��9�#����)5ޗB`A2�;���͵=�P����ƿuygw(�$��[�_]�^� �y�� ���o�e�~�P�|�w�jecZ��
��Q&�q�ךo�ϯ0�k5�V�rl0G+#�������_Լo��,�f�+*-u<跶 x�/Y��(��n�ޅ\�z� �F�۵a��W��^�Nw�z/��J����v	���
��������ا���% ���-hwܚ������o�����e����aLH�	!/F�c��;��ԗ�}����)�4�f���
3tvJH&j�|c3uC~	?E��F`3m���/�?�`�u����o��	@M�X9x�#��8�"_-�[�أlŵ�^�j��>/�-C�F�m�3X��Ȍ�fD
-� }��[f��.r��9��Q(�Zyi��¿_�3-&r{�0���-+��#���[�v� ��`��D�Uy����k#)�H-+�U��|���;hp�t{��7l��u��]����.��Aw��;ֻ���㜼��^�p�+75�3�����/��6
��@����e���s�D�0��6$����g�f��v��aj�+�1�:�{���زhf� ��1�]�)��\s�����a��sl�!N�O�/��1��u!�(��h�n�2u�*�v�#*HW�Sb\E���Ql��'�Pn�2�\���8�<�d��uGA?,�v�/k��nY���1��ϛ�Z�]��*�>���e~Y9��̮>�����8!��*�fk"���u�u�(��G�|J�z��;X�"�'A�p��)]�s]�};��6�v�©�ٯ||���?�mF�����(�g�wtG۪�&��TIZ����鑟���XQl���O��Vgɟ�1�9V� KA��KS��?�D�IVt��]��\\$E�kj�w�褢���Eh$d�������Q.�A�l%�g2��Vp�6J��j�	
��C���Bb¶M̪L#Ʀ�����:[ �Ʈ*ɓ��Wx����3���'Н�\d��O2#���ccv