XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����M�.��ka����[s�a���*�OA{`�<|wL��{\ [�ka��Ȓ��4��ͳqcF�~=��N?�!�b�:���V�>��h�����^F����B�%�*�:-���6�q���0G��������g����JI��'SCp�H1��W�ĥ������ǡIL�^���6@~F���,�������{��(p�M�VK�Ic ,4٨��:Q ϗ=@��lmL3y��;��ݹTG���e��f=c*3H���M��ɫ��NLCi.0���ٿX�r����!��|�4�������Y�_:8 �^X�D-d1 �[�
mD�3J e��	Q�=��Z�?5t�_��j=���A�R4�ҭ�Jzz��O���X*4�����x�~ʚ�劷������mb�䳳�/�]�N�ͬ�/�\F�Ŝ��O�=ȫ�I�b7�>����[T'5v��j������Vũ��;�Ӏ.����p��ޠ�����M�ħ|�$-r�ta�s��	�ׂ�7��ca}�Bm|`�sE�k+SZ֠�4�A;��BSs�x���݁@�GQֱ���Z��pb0��	�Ր"�a�dW?Ii�r�M�����y<����l@�Eu�ɵ�N��C��h%�#<R,�D�'v%�5�WYI��ۻ�s��.���DKGw� .��Iϝ�����sJ�s6:H`�PD�7���~fs�J^C��B�<Y���J&�IJ�{�ʩ��/|ЙD�)�Ep 鍗�߼Ң���W�Ed'�YP��LXlxVHYEB    1569     590&��c
��櫙�F��x~�2af�y���_�*1H����9ql�rHR��w�W[ڼ��C~#��#��u�Ğ�~חB̘Tmo�����ɬL>�z��~�bz�CM)��S7�[��ڋ[o&M�7�I�w����(6�>��_�wվv+�;�hi��o��Fk��Bp�7��Lﰐ9Sx��(Ξ�����ž���	���$*,��,j����YHu�?����1��H�+~	�O���O�3>��[{�����3{h'�ƥf�� �;Ԉg=D7dC i[�f6U�x��K��`�WSK�ݤ���Y}A/�;\��G�i#R�O9�g�G������hzd��[cR�z}�{��+.$�vv�~��'ꤍբB�~(ʡ�� ��җV���8�h1�E�1XΚ���!v�/��H�g;���S����L�{�?��u�S�R��R�~�����z��yfX��w1��b��V���B)���R��� Q�{nu�<n�n9�ɱ$n�t���s��nbz�X��{������v��,��Y9|�̖&R7��>��G��ہP\����F�3�O�jd!��[��8�҂���&iEX��a�@��Ձ
���4DK|	����^c�M�X���3!20�чe�4Ŋ:K�y�k�?������Px��V8ԨaL�z{f���6�N�����e>a��z�L��0�Y�L����1[_nO�.2{<�+�y�޸��wF��N4 ��_��l�I/����E#\֤p����;4V%�#֗�H�63�MZiD���3d�5J�yU?Y��9�\�����Д*5��$���J%�ʩ�.uX�
ǭ�(����xΰ������P5%�@��2��x�2l 9�����UG��p�'�|��W��:L���V!u���| @�/u���:2��|A�c��!�)��~%�����(��M�y��m�$�nՊ�)��]\Cw�4��w�iM)�57��Ͼ�oj(��J��2S�J��Q�s�Ĩ�d���M�]Ó�\����h�W��V�i��1��}�O�bz-&�0��T@l;\�6�K=���%��q�ht�0�qD�8�N�2�o�}���C4w�������W��������,��e��`mU�鰏�G~n����F����e�e�S��<Ȧg(�,��9�J�<\�0|�K���#�֗%�A3M��(r(���uX���[���N��)A.L�]l�McxJ�������?�/æN�xS�>/���Ivk8��X}"��f�W�I�A�6>X��o7x�"e�T�*\yעC��<��,}�#�OvP����o������a�β�s�铳$��Qt�*��6���Y��=�`g-�YT|!�6�[���3���K�k8�ꓽz}�h���pI�
I����