XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����U�:�1�$�a���z}���E���'�+ZC��	wO	I/��# ����9�@���4�=�����������a�rA�{�z�#eP2���Z�႐�����ۂZؽB2�hy���[���4���J�͕��%���������CM����xx�[C(��]���L8�s[-&�`2��	6���U�th�_4cwW�\ڐ�������6���u;�����	x��G�����TOq�8v������h8��ӎ�����#�6"�IUB?����6	j�&��C�.�|�4_�
���� LV/�W=E_S�Z���y�_��jϝ��P+T.�g/g-��~*v�N��T�2J $�Cӧu1�;k]�a��w�Zc�JZ�g!����j����yD:Do���Mj����4ޒ-�ޑ��Q"T�J���&M��d��ٿ7�k�V0�v����{���ا)�^)��\�]��˽��Q��(s�:�R�^��b�tT�L��N�����$�N��LQVd$��f>�D0����X�
�f�>����"b��ϛ�QE��� �� �F쯯���7]�`��ʐ��n��r�f�p������"�����F�*O�t(���n��,��3���B��eE�U#WCS�S��5�f�=�.ip&}��87��b��0z5�.	�\���8�ݦ���|ٳ��W�|}��z��62��꼭[0S�]���{��;�eħ���$.�%����Z]����⯴�m�����XlxVHYEB    6fc6     c30햞�ƥ���ʎd'0<S��/�|��=�j���	?�S:^{p�0cZ�p4�iiZ�
�b�xe22x�w{ �S�Q!l�٠`�u͙�6Ű��e���,�n��T󴹃��hVs,�jIy��Лz9���1���VӓLsʄ3Kn���Fy�.�Y}��
�E�ԛ8��A����'�-?�����`R���Ȋ��Z ��=����~�Ԥ��V}K�' �܈����U${��4���Q�)��״y�#��$���Z�,�`�Yw�0������#I�#���!<D�A�0��r���zepj�w��!?���m�6�3�"���c����*��y�.�YQi�R����(�����>�r-�Z��jR�*G*���F5��BئV��3�$��u�hI�%,隼5�jR�9*��:a���CW�n���2�X�+G2�*s>w��x��Y ��A��8�+����,��ԝ��2�)�b03q�fw�s����)��j��Q�h���Yw���Č[��Jl�ۢ�u�L����Cκ)���b�1���"M�:�UwԘZ.ԦFW\2�0L6%+i-�Ŵ���Yr�Z��&��ZI�%N��;X�B� oL%�p@�H���i,
���Yn �.=�{��͚��Qge��S�Wd`�۝j�'F�l�N��Hi%ҥ�� ���v=L�,J��u��Ū���)��1�9�r�n�����r���2�D9)ej@��{G�U��G�����-������a�w+'p������ Ig[�  NH��ُ^1B��mP�,�x|%_ļ�K�H����dY��!��<���Ox�Rb�ݞY޴S���pS����z�m�u�RP^{<��~���j����ttmF�
<���)�yU��������-�IӅ�8�kq��Tק�, 9*�2�Vc���2?3��c$����XDM����� Sf������aL�:�b?�T[�����Q�O��C�#~4AE�X?�`��F�H�^?{ ��d6c��T���o1���O��Sj$|���
>���W��b�q�/͑rEf�h�����J֗?��kv��x=#�;����߶8ޞ�c��4Q�C�?>���p�9.wa)v�9��ZI�̡���1��%�bA�.���M� 0�d�	-(p�.�l���f`�]�(r��@��&$�-v���Dǿ���r�NA�G��W�����>GSQ��m�i��8A��7�=��D��g��_u{�_�����7S��ȯ�K^��<"���k�Y�Ms��w����
b�)t��N�9&�O!��td���m٦?�)Y#�ǔ4 �w��rfc��G���e'�Sg��a�]I��h�0|�\ĮC�ư	866˛F�m+�Eu�0�o&p����.?�̴/��})�TЙ4k���P�t��z馅fUX�~���e�}F!]D�|�R�w���ځ���k���3��Њ���C��_Ori�.<B"�IO�"j�=w�R� �om𓆤ʊ�� @����V���J�Ps3�ڱߡHRl��m(�䱡KH"V
:3������?T�+���/eTP��_?��wpY�b�n��/A⏼�r|��7��V�;���83��*�@����_���d~^��p
��k��"���"����
P����S�c��=��i0�9�(T�_m�B=�d8DG��ъ����i_�b�9��(�G�r���~��j��wjt�8�,y
s��C0}9�P`4,�����߭����&��Go"�-�*�<+��3����Xj����)+♠c�M�������"�TS%�/0��^�f�f���E�%5a-�<���q��Gr���?�[�j��}�ᤶ�c���.��Ԉ�O�g�^�V}���y�*ќv�װ���H�*�G:Ew�(�k.�m�+i[
O��-��Ս��W�H�f`�Q<��Sg�|YT��PЫP|�{.�L�U��Ӓ�OH�@��� ,�64 ����n�*����@��$���x`,�8xt�wm��=����V�8-�[*B]�7��C�tY�=P+#2u��T�Qһ�{zB���A�)�F��������9��N��G��H��l]��-�yV����U��A���HXE	��i���r��DE.x��L���*q��x
k�����,�6��|7����^��X4+�j@��O�tَ
<Z4͓��bY��;�L�
�CG�����,z���%�;|�3v$;�2)~q6�D���exr��b�j8���*İ��`
xc��T���6sG����j��=޴��N|b�m*ܺ�]��e�����a�/~g�֘)Ĳ)� ���p��w⴨����~ ��S��a6�
�\~�B��)�?4W���)9����fGG���x�Lb�w�XC��xKR;i� �(�<�|r�#>E=3����eT�|ڞ������g_�_tVkz�A�E�0�x���T���{����af(���G�	ה�{V�`�Y(PH*e��iy?u���U�-\ѯ��)D0:cI*@�,h�O�p�Έ��{�Zy}�����;���`��3Kmdfz�FP+�6ٸD/�2��Ctd~��0Zg*w�`y�������y&���o�'�j���{�Kp4v��C�G�X��^�z��˒q���w%�3J\�\�:��㐘9,H���l��%��`�&�
��O
Ur��F��n+�f�U�va���a��s�VͶq{�}{�R��F�������H�Ws�SZ r�o��f����l(�xz�>��2�-�D�Mo���3�E1�oQ�N}�5�[!�܇�_hE����\��v���Ѯ@I��F�D ^������ӷ����E�%�(�%v��{d�2:��=o��,7��(��.��5\Å,8B�@�AP�Yh>�m�(&f���/^<GA$�Zc,�!�������,c��`��@�O>�	ȋ9�eɅ�.*�V�iU�VBԵ�[@4xS��Z�~l���Z��^m�N����s�� N���)����<��������ҁ���5�q������\��'�Ip�m