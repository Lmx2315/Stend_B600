XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��2��HM�!���0��:KJ?{ ��Y�1����K<��s*I��=U� �0NPT���F(�2 k:��%�[�G`_PE;n��0�dY'K��ty��M�a� �q솫e9K�mfD#a�x�q����h!"|E-J�KoJ�!�Cq;n���D�d��%B���ճ����ztʟ��{_��Q>��^Q�mu);<h���&Ra���Nx}Ny�bg��1OX���S��=[�B���an�ծ��]0��C0�G�4zY��c�j'=���րp�O]Մ��8��[�8A�%���K������F��ZѭUK���V��W��0ޯ�m)�T9��]D��j�c,a�T��'��CR39����~�08���M�+L�	R��1#�+NR�� ��Wm#Q؎IX@�F�8 u��~�ƾ9R�f���g�9��X�;�Me�j�y��DLŢ?�¡!,���4L��&�(��6��t���
�����X�U)W�����zhgUbH<u�R�͈�f���'��4�����k�?&��F�ή����U�r�� ��`h㈗xр���[�� )��NKD�_挺�߮�=��ڡO=���9]4���v���S�l�!�U������ɕ�-_�&-� |�w偨+�MН���L�w~�{�tV���袙��������:�G'�'��bR$��A,D�{�X	KC��B�)czZl�e&&-��x�7F����4P6�X�2OePb���7�	|tv����@�
�1��XlxVHYEB     686     2f0N㊟uE+]���W��[�����n���WSޙP����\�AO�;�`�m�wF��ؿ�zrI���F�r+OjE�?	@[��=HÆNS6n�:3��Q�õ��xh��(1$ۮ����(��#���66�۷9�,����g٭I�%�-��W������0���3nr�w�/0ҩ09���/�c�8��/� �Q�����l��+,i��BY��)�P�Z��G��k��P��M��4|�7˄g�Ų�|�E63낝�X4"V��e�6n E�j�_�h��:Ю1Q'lBW�0�B������\hN� s�l��t0z�!@S}B��hP!l�����^��gBC��̤��rrȤ��W1M<%���:��4jڌH����G���aa�H�X�s_�z�d��m�0UHNf�9��*�Q`j�wq�:���$�W�DD-�I�ھ�W��;%J��0�8RH'�U�G�1z^Ћ[H�}QDI����닑5!j��i�����s�q�{�	���{���Yd\� ;�Oq����Q�x:�כ�>�Y)�~+-��!��֍6��&�w	)_���q�h�&O�����A�G��f��Ƀ*G����~�(�x�c�^
A�gZq���s)v`�"C^C�,A-�$�2r̽c�@O�����Q`7��!I�G����.3��~OnF���%���YD��@<P [գa=V�y��p�� ��.$��|!a���i��,O�K׆k�(��