XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����������w�#�ݴn�ԅ�E0�	4T�2Jn�#���:��z}�x�m�N�È�d;�_y���_X����l�M���o���״�d�̃]�""�LE���V�m��=1��P� ۡ�^{v��%��P�k�~��ĜS8C"2�迎//�W�%�K_ s,8�?��+	�(]���! �.�dC����5�>Ҁ�h�r`j0į���Nl��i�}�R� , f�0�a����:gE�g�!�	l���<Ͳ����5a�m
�ٶ������tl�S��N��%V�b��Qr�HU��Ʌ�8�z���p5��y:��u3�)�;B_���oi^~�V�X[��PCo�C�U
��:`��&���-G���d��]"���G���f��С3L�<�HE����n��R&���t��
�m����h��">��U0���hO��C����%����y���ʙ��w�h��g i&4���׹8��]*:[�$����7?U�P���7�2V�����J!XJ4�"U>��$����|[n������՟��})e����q�,~b}��{��@��`F��Y��L��	�,n�*��B0?�$7�9�Cs,�Y��u������U��~�`�'><���W����c�Q����.K�y�nQԍaO����G�({�QF������ >�1��f]���ܘ����!���`�n����W�zXΥR��0/{:���������P�=H4�#���R�e��0To[XlxVHYEB    4a09     920��)�����ԅ�"l��Ε���c�k��ތ�S��_.�����B�*~�ֹcl_�����RH$�P)gT�=���T�'@`o~�x��:37����Y�ӄ��?3X��t,�'��݀9<Fx&-Ȼ{pܲ���-GE!�H*��ͥ8�����U����X8�����6��8W��p���Z:hN�`zwn����W�t-��>�FԜ=���>Yq�/,��s���^]O���d�D�\��ݸ%�<Z ��61Z�8�J�����Gn��:�h���u���c����t�r��|�x
3W5��V�ћ"F�²�2�����Ȟ�gr��Wmx�=�ޮu�iy��o��}L~m��-Z��
�l'!=��Ȑ����{/k�!�g/��o�9"�7,@����v��P�ޯ�L3��8�"UEsX�0�_x��Ʒk�Fy�Э�+�9HV�)�"�u�C��!�S�fq�*L��������H�������q�"G�?��KA�Q�R���J���<�!��o_=Κ��
�r���˟�Dv�W�}J�/C�
��zTQ��ʯ�v�KH��BF{���_P�RAg2`�s����?%ڎiB�^P�C��(�t�@��>�F�P,��c����K?1�j��c:J,��Ƴb�	���5�C�'���5&�(���}����9���?�X�lR|n+U�_��lr���yޜ�{��V(�ýK���>)�%��6���!�V�u=�,m�
��5^��α-�Ă��	^��:�<L>ײV�%�<퀜]����%�-��@�D�3:��5���Rl���η 2���������`܀���Q�q�㩮	�L�Ii�h�R�![%��'x],�%]�l�8��6�ٯQ�,�����6Q�<C��������Ŭ`,�L��ޅf��ݼ�^�^�YY��pr%-g�@J�WQ��WGA^�v{��؝k`�g�uPN#�i�t��e*X��#Ϣ{��7!����+�{�m��AJ�qj��W.偘p'n��� �t�������1�����!f��:��g`���yﱜ�B��d��������!4�����/����D���j��Ç�0=��7�r#�x؀؛�z`�#2�PN iƤ)����eA$5�qYnt��&Y�[��RӒ��u�r��z�g��	Y��(#5Y�&��j��@�eNmihVh����<��!��-�i�{f��Zaƿ!���}z7��z�l}�yw���#��,RhzP�xh��TR �<`� <t�X#�v�GTtYZ4�iү��Y�
@U>�#˻�1��JX�q�)�w��&|D;�ҫQ�s�Z��k+�0�G��J�p��0��e��9�	�5��/�<��r9���~�8���0c�Qa���xۧ�n	��N�mxͳ�FY����cS�6�A3�c��6/�B�N��}�������SJ�!{`Qt���@�d�B�,Ӝ F�ݲ)9������8O�N�Ē�e�����<��#�;6�i���]�	�A�(T�܀�'gZ��J��j1񭥎�wBb�uw����FF3ŵ����[�C*#�HQ}�-F�ms_����
�
š\�):bՍ@s��i��,��Üb|�3�x���K#�ZD�J��֭o�[^L��u�_w�C	�ӔM"dj����k\����)�_f�a�x�S��R.�n������&�&)�%U��7_6J(8�1��>r+H���1����}B�/�sRN;k�W٢�ӐR��V�!�|������/�,W���Z��M�d�z|J&U�$܅ �W����qd�`���d�p�"sK9f?�EQ?�Nv�r�;WU��ʉ��u�aN����l�\;�1�d�&FU1��S�]
Ҷ�@[���`r!�k�pa�C'N.!(SeJ�h�Q
��I���Q���oҦ@S���E���g-�3 G�`%��/���E6`�΃��j�O��_�R�<R"��"�3<���P��Q�(�l���מ5E��1(yQ��h����7�?�o[�,�Y-C�Gg}�PQ�o�_�;�{��禈�I�\T}ْ.B7���Y��ߝ=���g�wb
������ٻT��}�T)n=���.h�9���0�"ĵ�c�)'癛Qer����I�f%��<�k��[��Ff7`��	��goȦ��C/�E���S�c?"30N�ȅ��Sx
vbβ����cA.���uA;��
��r��$� �����Ė푳݈���F���U|���&Y�ʿ3,1 7,sb�f��
v��v�n��}����ʴ8IX�