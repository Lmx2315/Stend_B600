XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����H,��������{����K���s��49K��qvf�֖�5m���UB'Øǧu���);r"���3��G�Zھ��������|���]��|�ǔ�/T8� ��ro-�9z�!���̵^&��n�0b;�D0NQ ��CR�h�K?-��_]���w�V���/,�M��I"v��H̀|:퟽��T����"S����.�&�نR�k"�랎�^V�_H���	*?�aj�`�.P�r��
۸#���,��{G��k�o��h�	�����T�����$v#�1R�Hͮ�m;�:*д�P�\�t��H��ş�������NvɈ"��܇q�~-!���,��K��P?�-�DB��0ws� ��;�$@�TJ�+1I�H8�N���� )�2|�r��2֌(�˟OQ0���Cb̊�*zU�j>��\����k˪'݌��Z	�A�6���҅��\�4�Һn��'���z�;�~�vڿ;��W�nZ��>�#��3%�Z@%&R���/��6������-�:M����+��rCmR)���,y0��C�� 9�d�8£�?���0�֩���]#���	[h-�A��H�8�Z��k\�b$\ʊ�����ŇyRX�fX�e;�auÆ2���B��ܨ�-�������SI��L=�d�h�y{��J�?	ߠgTL*M�w'��ӯ|�0�%���	P�W.���(��V�9|tro5�C|Ì�Ѧ��_��@��XlxVHYEB    6408     e20gHN rW�� <WHx�rY�I48M���j�3 &�;�^C���7�-����4�B�J�M�a�T�f����h����Ʈ�q��O��G�h����C�L�4��e��"tŠoAlp�t����>E�5J�~إ��ND�sDe����sʽ \��_����v)Z/��Q��4'{'�,���?�z��#V�x
@�-��.��XU�~����Mdp�[�����]�n�X�����~������y�2!�6#h�6�`(���u�)�g������+��kq�$��3�89������ʧv��%zCܲ�4:n��W��ߏ�@��> Ȫ��q�&y������-'�6W�U!-Gy�Rv������<%]�g�ӊ����K�!�i�q�B2�BI��V4_[��GdX;�&�T� ��pL,D��`�F�������%麪���������}_Kr�K"�1�
%d������f򣢺�`��`��E)L���^��������:�1Ί� ˘�qYQ/� �\��{˵A����w�Q�ְ�G*�@VOV-���K���x���u�s�̇������k��Rۏt�B�lm�=���K?�X�J��ft�A@U�-�8۞�����Wvw�tJ��nQ	yi	i�Qn��(!0?Pm�4���?���*����l�`7ڱ�(��r�ǩ�jt����-0#M1w�Q�<�>�K}��������G�OI
��s��&i�,n��"UjƩ%/��($P��j��$n"fث�v���ns���f����hf������5"��K:6%$��r]B-7��Z�4���v*5�0��rǒp#�C�T�E��#F8."��=��߯�u���pw����z�N^Mk\��z��2�~!x�g�큪��r�G�g1Z�t�h�<[����L͡�E��[�-
��A����f�lP�ڣ��f�l�����Ԡ��ׄbi��&��':+a6� e<��+�"\j�@o��姍Nג��2�6o��� �)��n��B``[;M��.-4e	�it[��b=^>p]k�������B4{��PT���e&��{�nm�z���niX�!I	��2܈wLp5�M��&�S X�"��죗2�0�7��Q�:PnM���vtzpϱ�OB�*�_���@�aޞ��c?�!�����_�v,;]����7��"�7Q�߉��́�A�m_���T�U�(OoG�ag
Dk��ʚ�PG�g۪����o"����" �v�'X�G?ER���C`T��Q�e??ؗ9��*�C����x?hUDk�X��;4,-�h���@�b��J��Q���})dΉ���|tFs��4�_(6�	 ��~��g�,��t*�#N�z��k*�jƏe�1H�IoN��H��g��l�Ͻ�����)�>|y�Z�&�`>���$Kթ��K�@<t������+�����*hR�R+����, 9!X2��*}�F��^�^}%�o�+�BE���r��W�B��2ڼ�B��1:+MSg� �E��dr=E)]vۀ�.5��~HA�1�2��yM��FLxCG��Y�%�_P.m��e�P'�ǃ�^�&�	����z��J��'���gs�g�[�iȁ}�C���``���h՞[��^�����R�/�W%o]u~�>����,�/{2���1�3��A�O,���i���#}U���'�6<�:ꅒ{{��AW�F�d�����
�I��.��SS犋����� �J"py�B>�%�W_���&G���.�T����$1 I�|�'�������P��:YBR�z)����8�%��Th����lz�_+(NT���}�8���t�kp��z�I:��E�CH�������r�n�U�#�H����u�R�vKl�/��@&�-)�����;�ҷN��)�~wnKP�����k���L+���Ig�$*b�e.Z�]R6��Z���:L(����2`�,U1����m�Q'�e���j�uT�чY����BP����6]Q�u��l^b:�>��h�6t��I�Fؓ)�,o�̈�lq����=g�/{�V�s���~�B[1u�*��4@$ҽfY!.` =��N�CE`AD��T�ls���:�\��)�v���'[7o��U|��pU����l;	p�F�CH�o���
+z�nh�qa���<|�q��zčv6=-�����h9.(�Z�11�f��F,x��U�ֿ̤�������J��i˜;�UsĦ�A[<�ڢwZ�O,]!%0�G�җ���쪷���at�e!X�Ջ0{�Uh����GP�ǈ� ���6`d.��S)f��XRK��FH����,{띗oR@'��1�gN�ߚ[@pA�, 	�-��|T)�]���8��Ϫw}�j���E�x�����&�ֆ����r�/H�H�F����i%��Ue8�.�+v�[�ݞcǹ����,K��->���ӗ��l
�!E\v)�Z�$����;[ �{�]w�>�ϐ�� n�N�/Rp��+��3�=Y�A��c�F��:䧓�ԗ�0+��c���ȰR��	k���H
t ��"�AU�ኅT:�5�y�ƧY4A��넋�����K�1��U�c����=��+���j�%.�����y�OJlȼrC&�A>. J�`��0�F�/����{�Q�˃�<��R��ྊ����/�+���o*�^�'	�4��j��˴v8�`���ɉ>������r��`��/r�w5�3 O�q�.�&�<��['@.��^�rD�"�2^{q�P�RX'1��A3��|ky�i?g��.���w��7M*��3y�Y��5�Z�R�(4��k[Lf�B�z�K��F��gP�EX��D}��������˓Tl��NEQ��~=�����` �p��	��w�a�٠{��	��j$��Qg��9�N+3�h�Q-� �h/�nj����RƬ�&�;�<t�Q���eI}i�J%�zq�����S\�@k��H�����^��M��޵�k_7���$7��9�AY��N#�,���0����,�V�,	<z#�p�'і;9��x����V���xd�]�~�V�2 �˟�*�2*ߝ���(|��ލ>�@%H7t&=T,�_�GӒk\��u�U���g+�1cy��_�A��m}��T�I>E�1B�����t��� ������C�R���S�������mK�j�����IG��a��^�\/�q�C[�:+��w3��zn��Έ�;��+�7c��=���[���wj���]�x��y���݆̶E�x��G#|��g��O� n��9�����\��g[�[��}��Úg7|l��
��[���^��-�\A����h��\�0n�$��ϣ�9��S�Cߛ���s!�LҜ�wއ��ۍ��:�v�,��:��S�=��h0�&K�=c�$3�Ь7\������{�f�dl���e���ꎄ-�L�khx%=��y�Eygn���i�h�FF��o\N�,0rݚv)2wF����(h�(�ڼ���Ӄ(�@�!pg�k�d�RϞ~G��