XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��޳�^�ݡ�Λ�iLa��gb?v��	<<���
��@i��d�:�w�	@j4]��/Z��&��xUG�	�]CE�f'xwa�����߆�L��<�e���6�#h8�:���-�̹ԃФ��,�Œ9)Paʐ]�;1���NN!ْ"e0 _e�y8M�G#�����3�;O�X�\SY!V���+Zmt�H@�WO�����g�AG1a�5�� ���a}��e}��.�cM�
����i�X�D8?G,R�BG�KŀH��$`�h� ��WK��Q?�7�e�9�x��Uu�Fs�����N_�����h�Č��AM��}O��0M	�G[�2
�j�bzIl�e���.�F֊HU�	[w��A�������L��e�f�U�?;�,�]yI�����(é�4vfR�X� r}N7��W-E��m�� _����P=ЎƝ������A,��n<�8����/�)@�J�T��u���m��U�d
lubן�S�n�9k�DR�KT�P2J-�v�r�=>�֝j����p�@�j��M�"G�s�����=2��1�p�G2��\v������Fj�e֐�Is���%�?�Q�j*�-��cG�;�57v�����:�Ъ���&<�d{
�R��& ����F�4�S�U���e��-�Q��|�&�@P�U�u�Fǀ���*���[�$�?�,��ѠX��l�C�%��YK�yS~}?2^R��cd����~rn�)e�c)�p�TL�XlxVHYEB    1b22     760W`w�4J��F�����N��yt�~�unl1���f�n��[]��W�>��&B$̟�-����#q�$���\��,\yD��~*��
;ǚd ;?����5�,k̄���E&⻇K͋��βQCG���p��v�@n�[�@�Ι��Ə���o\B�3T1���<}�LL����P�`1/�'���oi��1���fm�kT��D�pͻ� }g�x��[!���<��&k�����@���a����}#����LE]��dQ��/�\���#�j��r9��z8��L�'()����5��#�X���N�%�`ÁR�J�ؖ�_�4�*��}���c�Fq�\��@� DV�Ob���<���u㲨s��W����/�.��P
��t��/�1���O�0�G�K@�z!gT���mGx�+��ZrL� �n�����i��?12�3�Ѻ�]I=μ�F:ek��ː�w�(��p<G��{�Ӯ`���G=�0���<`T߭A04�B�q�o���E)�Z����7� �8u��B��e�ڍ�<�fkV�N�[���$ݱL��sr�Nk��Q\.b�L	A�Jk��MU\���Y�a��	h�g���?�L��H�^�F["#S�'�MYYs��Q{�T��n����~D�8���$�L�0y�ioƵ�{�����A��݊�{MMYQ�B>wۃ�6^�i��?�zVޡ�J�g�X-R��z����%�Ph�A�r/��j���n�i��]��R`��4@����ȥX��w��hS5�-��gM�X}�+wo�9��3�b�9h�,�y1�U٫=����0��S=��B�r,������qa��93�g�3g��Kӱ��C6�\j]e�ś�D��U�0�G+���l�r���=��}�˩#����_4�sh��i��u)E��Ԧ�Ef˕n�RP�h�~/��/b������"|m� �M����>�x&	�D�V��*.�wB��O)(����i��O��dt���I.�,3<��vrN��ד�lp����9����Ћ+2
'�y&>>���A�X�E�[����麕���o9�Yd�(7墾�.�`���p�37������4-�;��2ZA���Y�
R�*!#{���3wTP�E2�Cri�ⷘ�i�LZW�V��k.��o�*fc�僪5�`���}N�sƅ�%�9E���g�]���+�/s ��XwЕ�vp�9�cX��r��t�x��%,~K��m��f��]q�����bj�xRz�.�E�~p���X3�x�)�x�2��8��GX=��ǍS����$��CE-��u�m�0C����Th�{�º�<���4��;���/n�6t�ǽ�q!�.W�%�}N�Z��}��l�=D[�KX9����!�Ԝjȩ�=��{N�DA���qp����7�3ƠRA����,����ᨂ	[�Vj��c���[-v�R�q��bh�Qܼ(�\��]��5�sŨ��&���"�?�2<K�G_q+ �Z�V�F��/S#'��=�^�D��������D �w�����.��_��{��o���m���I��3.v��[���c8������V�0�:c�c��� ��IA��%?����E����/u,��T6<V���k;0%�e�[Y�+�3޼�K�z��HI��17�nMn�}�.�
�B`I�#u(���*���l���?�i�!l
R6��w>J���ܳ�	�+�n��mycϣ]p>����w ����[$�����څ�[%�$ɹ��f�d�VZ7?�~�k8�<ʣ����:��ɇ�YA'�D��+�����0O�y]�9&�4��Z��Ϡ��VU���������fV�P�\Rf���