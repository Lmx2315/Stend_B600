XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����(b�J�[}��Wa����K@kA�����'V?m
���PmYL�u.����(E�W�6�֩?}�9V��Jv4]"]F�R�Ԋn �2���~W񪿿r�	@ry�+J��' +1y	H� 9��Rjp@�y&]�W��u\Ⱥf# �2��.��jۭ�Vv�������p��𵑂O�xHA�^�Q�9-
2W8��V1{��.��	�������)EI�р��}g	��k'��E8V.X�L6ؼ	�Ǎ$>�W�;l3�l�u�%���es�/�1:J�E �J������JYY���2O�m����c�}�B�1{9&�5({�6RD
L���ۇs{8� 5���$���x�`��ц�N�i���P=�¯�(����%�Ĳ�]pm�8�25믱?�@���U��,�H~y��&��B�7���3�5���Ċ�	���cR�i6?��i(g��6Xv6��k��Y7er�~�C�}�=���������L�����f�i�}6!g��	�BC�I�ĄY�l$R���3W�U	r:3�s��5w�r�g���%��J
,ystBqj�)X��k}���cu*y4�I�7P�0Cw�<L4V��T㉋+��J�:�aV��1~M}�W{�?H��vB<�dт�p��뉨��_Љ�td5M���n���`wV�S�5�쪺�,fH�^�<)�>�<]f-3Gۡ����r�����ٛ�9�i�z�G��g��T��� �~0J`fU����F�* 9�xXlxVHYEB    282d     8f0�5���,�cp�H�xsx=X/��%N�����m\@�+��U¢��t���[־XAv���%���4���鏖a��p��!�ٿ��C3�W��5��E�&1 ��F{�I�U�4��[�2}iB�L��آ.����f��G�����"�ak�+��$=#d��Z�`�@don�  ��#=w��Y�BE�?V�)>+�(��*��ⷭ����^�j�)z���\�k��oH6��y�˰���䊔�]�> �z--Ov<�av���k�o������hщ�5Qp��������`ʪ�ZO����p�=�r�*�K���Γ
*s2F�ϵu����LO�0[�9�%���Alg�Y��I���	r����h��O�_���X+xh?6�ZU�iN���ʲxk��2c�F���G�&�{� ;�iŌ��ɬk�V ��Z��"�&�l�� �g=1aҮ=A��o�,�s�(^�<H��{9����b��JVr�-����ݜ�s&z<�6�s��۪8m����qx#H[%{[��1���sPw`Ձ1ާ�ud�z�^���Q[�ɾ�T��_ִ��Nh�VܢR!�~]I�r<-q������z�������d�����$�6����W	6<e)�s	��"m�N�����G� 9��@v�͉�iM�3�i$�����7s-�7:��l�t���5�԰�W�L��R�g�r�����7�=�m-����ʆ
}LWqNC����m�1���<�#�����5R�a�����s�Ir�d-�Ԃ��S�m�<Lb^Qy�=���V��~R07ѥ@ͳ*,{�p�z���'%e]�m���Ԝ�}����v�����j���!x�.hY�!a��:K�����!�ӌ�;Xm6i�zc*��>$�������Vc��o�)���ov���mD,�[�R���߽��Y'��`ͯ� b�;�q��Rq�E:*�`�.ɏ�
�Ȧ��@���|�JI:2�F���-o�,�<�k����K�!����W�)0Pl�߼�(�ާS�=�, C���a��SΡE��Zw[��Y���%������h�L5�y�_�|���6��;����Ό5)6�!��
�6�b�r+%wC�F�7ٻ��<�I1�Q�rU�v�0u���?��ta�9%0����H'6|c�.�x��	�K�yD�yP�u_=?�QP'���|��n��eAa���-��0�ѯ��	@
���M*P>����#�3��/�Z��0+�_/r��oX��yނ[�
�Z� �:i&J�~��cB������L`d��?�����}��Q�5X�Lt�Ͳr4Y:�׭��٣C!���:�*�*yh�9����!�g��� [�В~J*%����C1�
�~A.�o���>�)���ځ���na����ݢE�N��$5,�%8��񐞊�e��Z�*��&���ő��R�����t����4��FF�K�䞳��C�KH[H�fS�$�2W�ת�Cp}��G*�2kǢ�b���p�C���x�eI���D���m��$a�6ݑK��Gt��A���mW��햰�|Nl��ㅟ2��D�H��M���:��g��#�+AG�ةd�H��7���!ԏ�$;`������-y�@�PA��,��߬���	�c>���G����uq~�_ ��;�1)JD�X���M���� �����ɪ�Pܕ/Mz?*<NƦH�~��}=ֻ��g����8RE����>�͖͍7v���:��S6V�.����B�%����+&�tb](7�*����2&j�4��䢳ⱡv�)�M]��/r������^��L9AbP9��y�U��� hb��,�9VY���?7����缨��>�-%�c��|Tf���T����	9-��j�0�_�ͻ��o~_T��%~��`˵έ�X4^G�0��<�/�v�9]1|i���2�e� +jJS��/f�U�"�%�"'ug#��I�W�#��!0���U�xt�HYs�]�TQO)7�vp�4̫�F��Nڇi}��|�Gl<����	��?�C�������4&BEQ�!3�� j�VOT�(3��S8u{ZY����:y�]0��X�5����s�b�@��jL�W$��M�ؕL!�;��4κ�x�kF���LA%'��I�	,.k����W��$����{��J�aT�l�&Կ�"���\�����tչ��x�