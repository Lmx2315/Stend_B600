XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��YD0�4��B���q�N_�ND#������R��R����D�}��ӈ����?"nO32>�:]
U����d��/cǞ�֖�
���j��0�>��A�zU2N)���v�,ub2�U�0�/��w������Co��I��􆔐%�g�zh�:Kah&�0��	)���B�)ZQ@��[��L�1��8�9$fl�O@ss:f�Ŗ��q*�[i7��`A�n����h��IGj+\䉺�o6/��'_Qd%�&�{1�K1�e��6�_�@ݞ}�G�QR�鷛4@����e�s�ʋ�{�뉵�ϰMj�	�@�GK=���O�{b14���!�Nz�1ۜVAJ��1<6�o� ["]����l�b��^t��&��2K��$� 	��{�u9�kG��$$ʀ���xg����F�t#���-����#��HF4��J:6ASȐ�uqh֑���<b��D=�<0!����z��t.�f���η�=̷��Ѕ�Z|^�tQR��O%|��?h
��s3�x��JyJ�;]�74/�0*K�{��f���oc�K�ǐ�;���r� �F.�����	8��w�lB�"|d���n�uU��I�\�;bj�����fƞ��]��yWN��ݛH~h�(�iدhy!�f���!Ѐ[��PU��=DFuN���,���G�Pz7�����[��8b��\D�f�� ��z�y���7�+���`�W������,�iȰS]K���f��?=�uAo:�d���W�W�XlxVHYEB    166e     4004�V8,�z|E�>�6���x�����"��P�=�"~L���%k��uc��Pq
��X.K��o����V�����>�9�蕣�D� ��]��f�ϕ�*ϑ�
�Gj<�O�m�6r�^�e������z猽�����EʾPA4�0l� �[��#����H��D�͈yÇTs���G��\x�~�/ƨ���$�V ��CJ� �"�T �[7��3?�u@����]�U���_�5'?�*��,�+����B�eP��5����>&akJ�.l�1���a���;�k٨��� ٚ�[������j���O��z����姙���7)y���\��M��c��h��I���^�XQ�~c����3]DS��9=5/�;o�-�LSw�	̮ag�D��ֿ� �g't�?M]o��nl�+�p{��U�$`TiD�����w�oLZ1t���=?[�v�j����z���~$r� eN�ţ�^��B�@z]1h�b�&%92�F���:�8�� ��3�P����'�$6-��	�1>_}K�>4~�7�"a3
?,Q�g��t�s/����T9(]XR��]�׽�0�e���<�D=��4I��#_p��S��>"��p2Vŧ���;UuneR����[_*�e>��5�uo�g�YG�T@Ɗ@
?3b�����P����)+�i�� ���8]͘(49�n/������w�o.�2#�����y����/ =���HP������G�﯆<Cc_R����;D�o"^µ�,<��3���!$�a�a��*�W'y[����{��3%�#�,�G��-b��n#J̊���>�K3 ��Cd��U�j��;h���7}z��Y&t���oy�I�m��5�^�bE��ZeH�����j��XVɚ��;u�>������`��J�:M#�����vC��_��f���3�ǣ�x\���~�rlc�x�W������'e�Y<\#1Pia��h��W��Τ/