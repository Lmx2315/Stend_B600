XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����s�z�G�ʫ(|���2�;9�oP�#z�׾�
l5�ח�)9$q����*1�������m�L+-~�^��d伆B{;�`HCl����~Z��`��cD�uf������s�<�T[��$��>���t�"�w�*z����/�T8L��}l�PO�� bVr�`Ԩ�����zx2Q4:_�x�l3{�ZD�[�-7jp��]�<h�96-���wZUk؁ZF]z'�K*/��������T��z�
�� Bd,O��{�[y�,�:q��ɇ�-'�_x�A&��D�t.�aL����O�g��Q]:Jd�a�����������9��N�� ���<�U���E�&\���� ����א��B|J� 0�[����5�:x�ף��8����s�g$�<<���0���5
�W˒�To���&���X�kZ$�������7|=���E�,>��q�~$<\�w_X�4^d��������;z�$U6�ꂀOp��P\�Z>�,�r���:������p
��%��qp��W�@:��`��C_F��,�ŷ��>'�ɠ�gk��?0�X߲�РY��5svY
�^Mn]����𣑀Ml��%��c�N�I�&�uB^��
H\Zd�����(7�����3fG�v�(���{�lΜ�L�9nr�Z6��,����+���7���A�^�̀��G��Z,SO�r�e�9O_��]q-���l�BEF,�e2���n�?��������
ǹ���Zb�+��P��9XlxVHYEB    4d93     cb0hH��T]�;F~�?BKye{�)&/��Iyq:�r�O�>
�A�o>�3�^,����t�ʾI�~Rȓ���jC�fnB��x�CO�þ�����3���69��.{I�i��N�q[k�z�:�=怄�U�%�25�U3��;s��,��r���vM�8�9y��"�xP�������qqF��/��L�	�/�1�f@���iVq5z!4챔u�����+L�x'�(����@��$�"�ta�H��|!3v����O�ZO��w�G���$��q������q�b�ڈ������0��~�2���r#:�|4�v�4�[ɿ/$%�o.-T�jޛ��Pn�v_���cP��U{�ܮ�b*9B]��м�^�^�^������t�h�@})%T�ːƟ�
��0���a� 
�x�nt&�I!�cc�O�_'����o?�P���l&�Y�hTXtT�:�@�ONV�r��F^�<�E X��0�{h�G��P���X3ePFI�e*���&�| ��Ͱ�<��[������汜x�e��8B��+��>�����!�z-�#�)-L��~�&�h6]���[.z�#0
�Fl �����1�uqڢH�\�SNU�TS�R�^������H�X_��hк�T��_l���YVoX}uK��@pD�ܰM�����uTj(�VIG�� �N�� �ʬ6��&Ĩ*E<���0	��l�Rle(���7�I�p�D�m�~��~�A 8�K?(1�T斚>��z�hp�1Q.O���B��t?P�+yc�	�&{�ٞB�;�����in ڞ\G����拠�%�9�Jy��b����e����R?Fd��0�ЀgD}�*w^��hX����< mנq�0B@����%��Q���^w�G�ח��$�-�~���si�[g�$\����c(,�����:��]�~�
�]���~��kP��lac�_RM/SJuf�Ы�*���=�S|�j4���zp��[%�;U�s]�(H�����8�6�s����r�[)W���a�J�,�+��h�}��������B�"^�Lꄞ�^s��+��=K
ڮ�V�b5�|b{s��{L���3��
�
��t��-���[�<$&Q�������Gwߵ�$��N��è�1�;���^Q)��@Sz@
��f�s��3�Ο+�@D�*ƗW���)5.�!�`��~���k*���1����r�'I5�h~ܔ��<F�	�^f�\��a��8f�O�B�Z����m�0D��� ���0ik3�])��h��v�8��Eܺ7��\5�k��ŭ��0�͗DFU� �e�9:�
"m�Ҧ�����?B2��|�t鑊�0���M�l:�x>1�FCGz3���e,
)�ϯ_M�uԒ�|"]�P'��ǷI�*ba�x�^W��
���Q��]q�ۂb9�Ϩ{1�^3(��Ɯf��D��!#V�
��h�Yc]ۤ�k?�<UFZ%&%y��\��Y{���;@�O���D��;r}���|�t��
PY�ކ{n�&��C�_K��m�p	V丞��*����/R���� E�ش���`�T�A/�VDY�GFA4=�-X�&l��@짻T���r��Ʋ}Mc4�aj��w�>D�!�p��{1ͧ��$T��$Stz��2���k�N��0foø�jH3�l3�@NT�e}Ne�0����� $���N��QTU�)���8�K;I��):�H�� #'���-_�:afҊ�g����V�J}Υe\C@������To1��[�E%����\ؒW����`��m�(!W
+m����`W�z�M��������l(k���;��D�D���i��~�aZ׎��-������JHị�HG��Qk� �r�}7P��!R��]y��^��o�e�Xg�����+K:Ϳc ��-�h5F|Q��%V4eֶ^���F�>�.����7!Pk\X�ڴ��m�N��HFY],�O1V�+`�%����p�T3�Yy��	]�$46	�����P� �̗�m�Ess�=fFc�/'?_�}v�c��7�R�:��6��<�w�_�ր��tz����3 �����?������1��^�����|��G�
��n]Kx��K�,��e���i|+��S�'��L�V�0SM�@-�k[�-g�w_
�Y�5N�}����;���W2��\���`��YHW���%`�CC,úo��	�*�"(އtLS�j;��=Rb��/P��u���w�k7Y:v�З�Y���h[�D�-e���Q�H�1�t�@M��Ie�IL$��׉��q�w����)Q��~���Sz\�0�Uژօ@b�dvv��L^pg���s�ȷ%'^q1[���"r�Ʒ=s���9֩5դ ��H�tNy�R��j��PJ:�I�ȋ<��%-\�>���i�����hN��>F�
�H�" ���V���9cM���v�!���X�98��9������[bm�N����9/�&*�I8��������<�'�(���E{$������Ʒ
u���
��E�{�/��&����|��/d�]��շ�^��4z�'PJ���<<:�Ȁ���x"�������d��t���\�ǜ4���`�����d�6Uߟ/H���D5��`¯2{�t�	7r��&���b�9��xג����j ������`��E�]Pf�����~�o���I��W�u.-g"�E�1���W@���ʳ+��a:ƃX�h���Kz�,P�BL4}�ۓqɳY'���	�Evr5�g.9����dߎ����Z�&��> �kO5 DI|���n��#�C�|����"�Z��ub�S��3���D��W�^/�v�|�z|��G��8X���f���y�
�l�,��9f� �)����r56�F����Te�W�ɩ^�j���D�C'�,V�"�~����C����m�pK;�,#���8ښ+3�!��]YÕ$Z4�oe{�~���a�|��:q�4��	dk���{� �.��cs�҄�/��Wܔ��R�6�$[(�x}�0�̋�O�u�N�+9���'ڈ '��U��yVR�3�R��˫
-��
��OB8Q���>�E�@�H����	s��GA�j�E^�k�*E�sK��˄SB|EGt�p�8�cinH��9J�N�������P:;�e`V^�w