XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��<�M}Q�e�u�S2Qm��j,}�J�(����L������Fv��RK���m3�g����M���mGf2���>e����`W�\QYXi�Zx�c�FD��N�u�=�φC���z@�S�Q��h[r'p+�{��R#Ű`T�*ho��ŭ�A�b�VQ�$~��j;�5j�@z܅��*Z�l��]�����1*KD�x���煉H�Φ�ģ^q��?n�q� �ZV� �E:pa)q�,&xN�D����dT>��C���+��_6�it�y(b��N�|�r��ڸɫ?�� 6M}�����]q��$Ӥ�T�u9�/�	��3䬒;G���Zv8���ni�6\J��.(���T#%*�����"��,��/���%
�3�C�!Y�A_���a˱X|_1�fZ5*-)�A�/������Ĩ��2��p�� ���,X{���@3J����4��?QJp���t������zf1+��n��/n�B��#�$��[׿4~髚�s��$i�I}��AG��U3*M�I��V��!s���̹N��$��S -=�Am���.l���I ��� �fڽv�V
<��L%ڌwvڠuP��M������rt���cJÂ2>uM�_K9l�Ir��3����*_<-Щ����j����O��4�EsH�ZS���ܴT.�p�nq�j8[���g>P'n��*1�LZ��]��޹p�be(Z]��{��Py�b��3Zm"uLp�3<ШZ������n���.�$XlxVHYEB    1cf8     790���"�]�5��������gQ�e73N�Y[j���7X�n�%cé_Wď��ͩte�L�y�mD-�ԔG�~���{q[� 9����8����V�L`_)@�8_�:h)�&GtL&�J9���ːm3E�o	1U���	Kk���b�|�uE�,@��.8���P���*�]%�y�l�^�;�f�i�s�f��v�p��!B
��������F���Iv�$���~%C��!F:Z�P�V2��of���Ӕ�(% ۊ��U��8ɱ8�J*��,hl���M�bh8�X���������Ff��K�J�l/�(Ƴ���h.h�	Ðj��ě� Y�FI>o���f<xDO��|Z��i���~�0�R,�jW�nW����-��#�3�6�R�o7⠷ ��vNn��E���`�Z���	-<ǎ��+W��ҏIׅ�s�=�S/���5���Z��< �
�a�ۿV6)Gt�ls���ۤX�9̠fl��"U�4�Æ.�q 6Z��;r�U�3r�?���#��vȟF�������#P���N[b��{f����U\%����&|vuA�?Q��%ăܲf����<��h�`���q�z�
E�ʭ�L�𮘀�E����&�����7U�J�"����{)�x�n��N�q�y�#�d~��g��
���#`�Gf���+�h��/�wXE��A��RH7,$4 ��Ec��߳���[��
��݀�cZ~���-�+�� k	�!Q�?�Da7��]x&Di ���Yd� ��V�G�x�Ȉi`iR�������b��rW�iE�|h��a	��g`$����U\�T"sM0*������D~�����2��Z�A���K(�Zb�Л}����a֎�-����{ޅjczާ��a{��T�#BL��Uq�q������t����~�蝈��`�Y�N�rB@h,�?҆w��k��)�S��`�K���0^�臟Zt&���(��k�,Z����(�M�	6dׇ�(�����X��/��0��_�(����}���-�sI���W�d��p�x'����;i)\�F?b@cw�xu깩A���hA����cF� ohKi�BHK�IJ��!�Vl�܆z�Gz_F9nkYc\�؍��,�*Hx�Dp�k�Su�ɬ�&���*6��$�!��<�B�)hw��.2Y鑖����F����w�Vؓd���?afϥ�e�-��!I���
Y���f�AH�h��&��1�q��5�����e��U�zh�w_�Cpy�HW�h>�Lr�2(�P�s"���1S's���>3.Z+�P5X�l^n��w�in��P���Ŧ�
F�O۸� 4!P�bM=��I�K�Q-dUk}�_R��9���EŜ�L)5�����b̗��K�vE�r�
NByU�f������u��[�i70hTg^J�:cpK��׾jJᛝ`=���HSB�<8(���Lr��P�I�:|����B��T��}�|������F��x�b�7RNrqT��/o��EG��q��A]�O�٘�1KxM0�fxF��F����5��M��r5�Rq���������W��/���h
�H,*��`�O�~B�d�a�Ԫ��<?#��R��Gep��t��9��(��?K�!��j���"�g}>��]L�D��x̂�㢮b�qG)@�J㨅�K��[��'�]��㢣�� K 4"��uj3�y/�dP)`���U#�R'���jA���%������=t��"neT��N
�#e;=����KF��v�;�HL�g��2�18�9��yT����Ae�%��ٹ�F��i��a�#è�x��ֵ%(�V�8���f��$�S�օ�>������󿦎�� $,hmŌ��W{�G�TW�e~�O|�6��Fr_Fwڸ�6T�4�B