XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��yib�r-@������{f�U&�咫���:L�g���&�ʊy��G���R�x�[�N�WGh�_B~[j�~�Ǿ�6i��ȝ\������T��X����n���%B��e�ԍ�i^�>����0(*�X�;M̮ߨ���<�LC�s�+����*�:�`��f�P�J7�����ֺ�����oy�Me�FW9���+~��x�7�Ȍytѡ�BH�������mx�ߓ	��%L�~jڂ�O�85�N�	��H��lW�N#�d�I�h�h'�@F��1r'�L��QI�4�����7J�&O8����E���)�[�"#���a"[�{����2��,�W���H"``:�250�Z�Ͻ���7>J�Nf�%���WV,���S����e�����P�kG#��
��B��<�0�LtGm,�ۨNG�`C`}&kZجv#$�7BU�Oυ�oj�~⨑�~���ϵ�p��;��y8�Ecj:�wtA��\3_̜�?��u+ޢo��V�)n/	��������S�]�A�$�		״$à&��8Gw��p�c����K�>�5ǒ�&��Ig҅)-B��� �M�.AG�>FR��+S�	����Kiv�X{n�퀶�'֪�Ѿ�'*ū�݄
L�!W���-%:y��b�DaXg  ��S���ݮ&S4�����Cގ9Ú��&|f�Q�hE���N\��%{����{2lbW�nȆ�+�n���J�F�'%�k��RM�5�1�o���+/���b5XlxVHYEB    6d0a     be0��r=�x�NY���v�^Pu��Ll�ԱEV�Y1!�
��c  ���vV5�|+>�V[M��
g�$����-�6��X��I���?ů	���#��Vh"�ű�Eq�)jOư�(�������7A��̗���K�sܪ�~�M�:��Λ�ݾ�.��&�R �DٶaTى��ޥ1O_���aMy��Ev����+��wW��~����X ��)?ǹ@��)�5 �(������\d��N�<�����f�}���$PC3�E�g�b�-"W9ؕ;�3�s��>��KW�H���=&q�k������Iҗ�)g;;����oF��~�Á��j!c��7��}Z���i�uO��2��z���w�*�
s#P��s��OxAϾX���OC��?3g�<�b���!0�R1�W+[�5��F����q���0/櫷j�ӗ�G�0k�]:�}��ޗD�%����Qɮ���J��-u�a�[��4Q����n��7�6�¥��f�Te��|`>}er���pK�&�U����jP�����PfWn����T5���,�0���61��s3�L�J|�%H$�%*N��D���|[' 4�q���qV���^
F/6���V)z�io�����8�e���?�����4���\�V�!���H�6�Ҡ$�FTm����u�G���Q5{�A�<��zhq��i��9�ˠ��@ԏ]K���	��	=��Vm	�C���/!�%`P�ߡ7����7�d>�������,�޲:�1 ������:��:w#�F��B�C��?�O�w�n��V��~~�B�.���=̍ �4��H!��e)=NQ Q[v�YQq �P�F�*�/�~g��}7<w��h����e4U�I�<)�����Pd�g���E��y�I�����F���.\�8 �kYԄ�l��Pa	&�]��m��U��@xv<b��7$sR;�	d��Q����̷T���Z)��C���������3�Y���d�Qt�2E�5�]8��g�B,�`�b)�A�2�ϱZ$W$A� �փ�yb�����z����g(&;����v[��h�ym��m]Qv<���T)Ҟ�$�-�NP�.� ����F��E��ǒ�PƬY������RE�#-��-���m"X!-�&��υc:i�x���0���&-ћ;w�\��7�+"K\&z	�K����,Zg�T�V��ŝk�Bd�z}T��pR��m������*���~�.8ѭ+B]����e��v�0�`�CiM� ���#�XjSX�;������wQ��r��$�O9#Q]����D��}AKz����MoI$dJv��YޞEl�yC���'Wi?�a��!�M>�Љ����H1l���y]�H9f�&;��m�e����c9l]c���[�(��TeT�����@���u�	�<=����������� 5s�ED����hA�&��n8{Ԭ�H�'�x�A�N�u�.pǏ��:MC�Ù0ef28��e�=�����gc�}�(&g�2���'^4���^�>Sj$3���+�����9,y���N�,>�܂f�g^�Whi�ˎ
��i���$ͦ��\���2�����e>Zd1�*��f�E�����+��z~?�1�u�z8���	�p��_�]!�Ӌ�q�k'C2�}���N���9X�k/3��f�zW���h�*ĥ��3#������i9��$��c���:� 	�|{�%�̇M
��b�IY�a�c��|jK�����8��۳���ܹ^�x �9�|�.���u�&����3�o�7)�i~�g��p�r�>�L2@;�Zxղ�JGE�ز�	�I�0��1;�SJ��{��5����>�$��>�a��<�h��R�MJ,�ӹZ�G��v65��ݐ�4�.Cs�\�߯4L�3�g�n(��W�:k1��l����0j�V_?�pd�Q�˦����R�`M��P>��0��d�Z��=��j��x�	��"��l@�_��:�n�;B���ݤ�3m���1v�q+>��[4�Ѧ~���&u�]DHf-s�ه�ڎ�ɶKm��t�#�e.�M��X-x?�34�HdʡT����8EL���Jp�ԛ�8���܏��I�y��}G������ah5������Vcb��Q��͐cG��9a��I�G3��@F��ks�<!�拾���3E�����f�Q��)	T?G�gK�{>�1 e�[4�dl�S(��o35��W��\��B+�j�����M:�a�q|��zչ+���~ ������2��$�\���������ݓ�L9`W[5���,��Bu�\��y�$m��ݸ����7�YR}��
��c>���FG6���Ǝs�ܷ�N�� 0�����y�P(�@��7;`���$fb��,��M-׻X!iǝov:q"�"�w%UH��7�1�����%P_���J2��{��E�xe%�u��Y:߀~)э���&�4& \�4^&�PU�c��K!b�U'�92��s�`����K�(������.��k��IA��b;&�M�Ml����L�#��/e'���|4�e���3�G�)>d����+���zU"��u/P�e/�)D�y�^��]<R��fӻs�K>�+���A��^GI�o�%�a=�ҕ��֤Z����.f�u${!���Q�;�c�ʨ
�M���>^Y�Fg����0D�|�3t#]#���F��G� �f�T����)D��uh��k�%eK����DRx�c�x+��f�S�ᾥ^�`�[OI�h��l��"�Z<���*&8��+|ȴ�73!�e�.�S����ϡ'EW��Mo����g��(3����( @��A´�sh���iU���i���}�xe��O*�9��c��d� Rec��'=�Ɋ�k��W&�?���,���1��s�&!��щf����Z��k�yxm��V��QQ_��E�Er5{)�J