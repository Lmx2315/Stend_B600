XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����tk�����\��ΩlT��� 0jz&��s�BfjY �l�|�9��+w9puD��DH]ż��~I)Y�bw��5�b�,;�@���h�>�A�!~L`�Bηq1�>:+�V�2�!=> ը���ܢ]s���*)�*&���p�si�gm8�kV)�gU��q����i�� i�����/~G�~)V%�K��;D�f�m�'�����z�P�]D���6lidD��s����6���[�%��2�&��^��ޚ���"䉭��0�tP�ÔYW߹� �9ג��S?��B�őo|'�	�<�:��1��@�4���ƙ�|�l/Ṣ|����g�,���ԚV��&����X2%2a���ݖ�����r���o��LB�\~��<9�W��m��Gf�Ʈ��i*		4�>x��f-��x����<C�{��[����!}�
:`;��ܴzR�l�>��5�k�j��,Qh�l��x�*8���O�'�_ă��ś���n�q�|�XEvW�L@q�zq�
V��7h��fj���.�r@5n�������}�R!E����;�͋FV���&|S���q��H�y�'�蝑'$o�t啻�H��o�̓���k��k����S�S���;�N^�Ny��?-2H��+�*�["��������ǗL���916�e����R�0��ڔ�����@甠 ��T��^26���/M�N&xx �3��h�����9gC��P!'�d��`F��~ܘXlxVHYEB    3a1b     d40�ź�' Za/�t�D6<�wf�Fya4�4�/|:8:����u�;����1�PO���K� w�\I�k����.f!��0��v
"���9��~��IQ:i|��'CǤ�\��yPC�OV�vNIaT����h[!{�0���Ɋ&����s����ڌ�bqiZ�6��G�J��B�',�$����z|),šV�����mҮ�F̿<jG%"	P�C����� �m�A�͟�S<!������>}U�Y?)����9�jw�M�q��~�쪛y�����r0C��m�K�#3R2���O�x�D�ޓ>*.����ʎ�-�r%�'5+||��!3s��cw����.Ǜ�Ŗ���;[�\2�[`,"o��*��\ӈ�+�{s�Ǧ��]��O��@�w�����n��s-�����?�4!�U�'yϚ���P9<"��e�֮���u� 5�m^n	���w��q�L�V��g~{:U6�l�i_�R��M;�Sb������)���E��Ǚp<T������􅄧/�~A5d@VӶ}����P\�B�Q~Qm��\�?y|�'+#`s�褨��>���gy�##^�dTq��sx��EH�A@	8E�K	!��i���M��6N. �w�V`e�u�q�@�}��w8�߆A��@%8#������P�5]�b� ��2(���>6GϜfv�9�[@����aN�S��bMگ^F�DV]���*d����s�3�cZ$'y�5�_?���m�O5����˺��N����~���Pp�#���F�C�8�ݜ��%C�b�1��<W�0sF ��u�]�%��	R0�sf�V�N0�N��״���W�憏������
gG�[_�nJT�%�E����dW��!�\�=2%�����������Ru�w�{OB��+R[�͋��&�3<������S��S���Zy��70N���+v�n@yO�V�	[��H�pt/�����*1ę
�U�~�W_��//`�l4{�9Cn)Yw�G�M}�I�7�ȃy��gj��m%�@<p���)�uc�з�E�Å���W��1�k�!D�7&���;}��L���wבtD0�D��]Z|r%)E1�.����x���X5KL�נ�J�|�%ሃ$JgAaطo�ݙY��l��w#�A'{2QˉA���j]�cW�#���ap�L��vs����+Du��%�:��Q��.���	̓>m��h�N�s�v���V��]"��x�e$/m�9�-�5&��/�V ��#�
�6Qpn$D�m4k�������u.���V���?z�FN�'�I>�t��9o��_j���v 5�R�@��#�9~F���+Ef=`	��`�'��5K���{�N����7����h�%G��oW�J���;jΈ���mw��2�����h�DX�>7��~�!���(�:����ؤ��| ����=����-��Q�i��I�^%2mN��d+�C,��lb��P��f�M���k����d��������5�F#e*Ģu@�S�ў�
�~�Rp̀�ET|w������N��q�[�HX��Q��|0r��ӕ���>a�K�\]k]�(�r_5A�z�4h�(hI\x.�,Ǳ�����TK�BU�eN2%>á�P�.\v[,U�'[����9Z�����I�)�弃��ɋ�6��+0@cĿ�]e<[�������3x�YKK(Y��BB�L0�UX�w]=́_t��9���j,ƀ𑶌�ݞ�D��gk��TZצ����v�6bƛ�Y�f)�5���YRMtt>*�[�j�����6+c|Ʋ̿�./pI�؟� �|��+��:	��'�+L�\m�h�����"51������t�q:c ��۹O{�kq���a̋��џ�1C={���Ό�� S%��5S#��"d(����lC�s6���-Dn/ܫ�ڵC�o�?�k����ߗ&t$�}?� �Bn��QQ�hF���T�6�=69�U�=@oIRy�Na��� �;�՗�pk'��c%8j�T]�v���J��Q����$���žF���r^�����(pn/Pި��4t�-ޱf�Iu��"'8��͍�b��|���ʴ7�}�1~7*LJ.�1}>��d�g��Vɷ��f�3UmD0z�ٳ�F(�h�TQ��jT#���I����@p�;�\�Lu
���n+ݹө]
��%F�{`��#��IQ�9�%����!��_�B�+��Q��	�F�����{̙"�z��&���2�bt.��7��y�Qݿ�-�L~p�Ӷ�e���n��zL�6����?�{h�S�Å`Њ��~�<�]M:�ӡɜ���ײ��5Y$���ռ�
�̃X���ޗo���]�^��X%�Cxb���s���؀'���־o�Je����	gξ�Yv
��T�5C��:��;.��z�{S���a2�G>:�E,U�6����ʡ�(�*�O�yH��ȏ�E���O�z��/R}�O�H�А�e/h%W,��D'�%��]0��e�zN�ӳ_�4�#�?�6����``���8-\�U5����7�b��79=�m�&F�X��`�x�zd
t�WV��yѨ�1�n�T��X� c�Z������.Rf/��z��3����U��
�E�����M!�Pg�Ui�� W��g��ԑ�S����Ic��*��֪P��;���,��x�,�����E����G���C��DŠA���R_������Dđ�3Z5ꘋ����Ml=YM^����(8�Q\}�   �T�K�P��)ѭ�͋\�>U����C�t ���W�?
^!�|oE�?iP�:�H�'Q�,��D�1o��ЍX�3}̫�0й��"��2�.JA�tilԤR��d�|��FØw��kQ�)�{V!��<ԏa*$
]�
|*���)md���>E�qq�=y����˵�� �)-7RS��x]��>U�h�"����(w%�H8�R+�"�{.�ȟx�D&�Y+	Lk�$-AWgt`�:����LT��B1�p��
���4��Q-f�q�s7�y���5�!n"1�C:2�s��52��2g {�0`�߿}����E���i�#M �0u=>�>+�7i7L��JѰ�>N������;�r[�#��>#,8�_K���ɝU��o�RP �������%^\_�P�YVv\
sʎ榛�!f?����HX$Ҡ�껔F�rkf��~,���|� ��N���.�t����8����㘻w�V`����U%m0�+���''W|y?��	{�	B`6%@��B���F�0ײ����e�:���A�WH
s(P