XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���A\)N��(w�٧UfS�,��>
U��r�O(p�L0]R+�nċ)��#p��nFa���q��O򝻻�okL��锊�0�,����=��p9�x>)� ��Pcy�"��NdhX$�9U��.Z�#���i5@���`�M��n%ub�kt��J�e�����TM`T~��E��K)2z�
�M*&��m�!��ʺ	b#��ϖ�MD�hxL�y����I�k@@�rz{D.��W�V��빩R��lm�)�\)> om�A��p��k�qL�\���l�}�N$O7���>�g�i�bp�׎�t��K&����I�����i�����'�M ~$wd/+Z��*�Z���r}N�i-�c.�l�_�S ;�]~X�ր�3����w1��%��`����*U �?�$Kv�0�D,^��"w�&�Ŧ����VkK�6����Ͻ�?Nj��l���֨7W�G�����h�Ad�Vm2�+f�b���2�(�EV�3���[26S��[�cp�C��?�\�;��1�nb"U�Ϥ߄K�VU��d��C���R�X՚��3�V7�*���o��)��-%80�X2#��>*Nqǂ����fR��tK �����`m)�����m:�� g�t���pGw��a�ܕ�4�	���F���\�y���bs�x��;��[K�ָ|8n�"G^'s���VS�y�2X՚I�:�����3�r���ح�����g���"��=P��2]>�x�������~ω��XlxVHYEB    2864     8d076�3���F]���-o�k�+8�Y@A���0B�c����Gt=j��v7JK-�L�|��/|�;��>+\ម����R��-*�ʢ�/?܆�FG��J!���MB����G�7���[�&����%[Ե+���.���:TO�y��N�I{B �u&a��{4O-+,tyɐ�!$�D����l��y��J.����!Ez�1� �\��t� x�����K	K,^넴L�i���ä��]~Pq� ��Y;H��P*~5��-�M9����m	d�[��8����vޥ�&>�F���[TtR�j�??DU�$�], ^���}��:��x7��JvM���-�j6`�b�V(9Ht'ƲF�Q���ܳ4!����;�🂇�f#-i�� �y
��{!d>������7Zz�Q!'�k�� �����������Df���--���0�=�� �U&��b����R1s(P�]�/'v��#�"�L�(��� ���x����[�D�'9�D�O�A�u�4^Q*4��
�{)������e�b�^�u0G����jY����E�N�6Θ�/��sT׆��
������+W��z�h׎:��1^���C�w�x�nM]U�ػ�_�E'���l��oj�P��ӠD{@skz5�(id��AI �x�l̚i��ќy_Rz�Y�W�I�:b�1��Ÿ�I
�E}��j�i��4���_j�}n�t2/�~�����U&���E���I\I8q�`�`7s�)�"�֩G�>3H�lv6%-���ҿ�|�GA,AT�2��Ė1SS_�34쭲u�;{9�����i�9P�{��cx�=�z&��*�N��v�sy��</�?#X}�o/���8#
j�jiW���<G!O�yw��^���
~��ƀ��{�]̵�߽2D���s�2�g���OCMgKv(j��W�fk��\�M�J鉦��r��E����Ǎ�nT��g�E~�e��52�ؐ��n�����s�h�}�x�2f���/ݣ�;���)H4�
Q��K;��5����޾79�׆?�f8	_�Wh�N(گ`�ʆ�ҵ<(�����8�.;��ħ���	aG�Z����k�Z��^�ՔܾBݠ�<��`�� 1E�x-a�x�}A]�v+~��is�Y�(���+����j����@1
�ׂj��t`���No�8�(�s�1�ױhU�;��ӥ�&P�s'����L�
�<	��(�.���wj�!��#o\V��I���)���ٙ��`���
sZ]y����;C\K���t�W�����R��Hg	����f�<�d��Gh��'�y�Ub7�`�MpP���4i����ӿ�^��%��d�M�ƶ����v��T�g�eUOd��A��͞�47�y.,�GF��>�4�
���g��SAC��?\�zgq�7��j�s�Ѡ���+(Kگ�|*"3!�Ă` ��Rl].�Sr��*�؟M� w�P�y�¤�o�y-f�����SN�'CTǓ�ay�}��l�ҭ���������Ձ�Oĺn	WXQ$�,�P�dYC�V��d4�`%6[|�����,d��j���`o�و��h�F8�s}�0�.���^�-��k�:U��8�C�U�s�DR	��+,�q >`�f<��e���բ��Z�X�A˦Z�]�
Qv�^�+��54��R��Jv�_�;[:�NI��w�S�n��GxU�����)|9�}d��@I�y$%�Wʹj�.G-Q#ԅ��\��yN~8mms�����˻FZ��_1������{�� �   ��Vm� {�
$L)���Ir�/oŧa�|9�~X��z��<q�ko�C�lփ��l73w�Y��4� �ȼGg��yO��&o$j��sF&&���	F
2�gVfrRr2��
s���s�������ɯ�K{$��ؾ��!�Z��M��/�ke��P���:�Y��-vŨ>�S�ߙ��l3}!q����p�*�u��-��a�*&��e�"�(����n����n^�g����N����;Yi��	�4���+�R�Y�m�}oJ�<`��-{�����?����`���ٓ?Y �P����5���*��� �1�:u'�Qh�ȆJ(��>�1|.�݄tk'c�mS��@�Yo����$��	{��w!��*� @�`��g�O|r@!�Sl@x<&�3M譭�~����&�