XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��9����TPe���Y��*фv��9,z����P�k���Gi1�һ��{6P�7et-T�qt�����"��nfR�����?�������y����;����0עȃpW�������ۤ)��!HB��$�o�i:onoc�Y!]7���x1]>�6�j�d�����.��nI�Ҏb5��]�(��k�v��|�>b�����(�	S�9Y��$~�Wi�1|�Qa;eF�H�N:��b�f٠8@z���C~T�	I`�І�(¤϶R�$S�@�9a�+7�&�^g�[��"7��ߦ������qk^�w+�z6׻�������:GySQ�~u�Z�B`cqcj��K�7��g��nxx���~��}�b���ׯ�6���$�������{��օ(I��a X�4p��/���	���̱:R4��'�~�L֟᣶G�LͧO��k�ņ��oÌ�`����`XW�ԯ�c�έC�H�_��Z�����ry���n�uxDOA�u�n��u�+�y�|��l�\�^t}�%#^gl�dh�X8��ŬI�[����_o��h�Wk�(�6�@������-�W&)��d���X���k��3*�����5��<>��g� ��>f�tk�X�~�%EpH<�0hC\,��p3٣R.Wyx����`�0��,�(},j��'ojkG��~ ���2���A��\�hDw�:�/���l���_O��J³���A�:������e炔�^劜pR|�6EN�XlxVHYEB     b7b     470��m�����3�9&�~��L�q�T�"5]�K��s���ߧiF�SV��=�����C�}��M�����X��GZX|����ԀVT�A���v2�o�������7@X���)�������Ã6�	��w���p1���I~��4���������]�%����P����O����E}6D��7\2�$�1k�A���M�E!b'~Y�l�Z.ƆH���$r�� TqٲQ?�xsT���x&�1�`�%���5�P�
�d>��o�s���Bǝ��~���nFk-j}��@5�q�x��1�W�|�{�I��A�nfG�4��>Rc�,|�fKb[�MFD�Et�gi����~˭L~�w��΍�a�4��$�Λ�.���9�X�JҨBE�8U�^3���v���EZ{d�j~g�C#N�����̊�_�t��q��z~+9�慠y��er���2[����Un�5��6,k|�8�a����g8��� S�4F	��zQ��K]��/����?1���w���<���ɳkUa��AEh��_���^)�a3@啷5����?��e�ϩVt�p}V�~/o�_Y�bM P��	J��k��l�f�ӹ.Pgr���Z�#N�N���
�%���*1F��W3�*�,�;������mu��&\�ސ�_����1*R�rA�x��O�:E#�%�G:�i���Ԭ�@�^�II��$���WTP)�7[���҈&~� :�ހK��#)�+�]�җ&��K Iy�Gp���vh�XU�_�lW�ۑn��:��ݶ<��bf�/��ɛv
�q��=qpw���5 �����1Q�Kk)�S�}�J�����F�0Y�;�;�۳I�Ag�5�4T8|���B��y&�B��^��|��;%���w1��/����$�	�n���eH ��u�n��Æc6y/	�w�rrl;N�t�e9���r6ЈBi��9��j��)��`N��7�����u;�N���Ն�=��䮖��|�J
����O5=L���3�ǿ0e
�Ok��y�pK�z#�R�ɡN'�Փ��|;lY�3�����jHIO켛r�1Ŋ�eS�ǋ�^���9-�Q-�:wD�>rƵXn~�'{����