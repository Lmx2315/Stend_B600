XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���%rgީb`B�ɢ��I`H\3lb� (�I�w���F�|8'�)z� f;�P��&)�Y�|T?���E��g{��)y ����+�����0ug(�/r�E?0�/5��ٗ��0���0Z?���@�{w����W�Ǽsu��_b���8j�I=|��9Bk�d�k�t�C���j���^�y��apvϙ�O�q��2?+ �}��\΋�L>��]NBq�@���8ظ��6>�=F�{Eu����<q�~�5蒷���q��!;w�B�&B�f�(��`�'�Ѵ;uk"�3��!";=�5'Zg&]�K���J�5O��UZD5^)x|��̰��̱x�� ��Ƴ�UH�0�ToM�\�3�WW�=Q,�:��6��?BR�xO�v�{�QxƖMܿh���,��;&���-���O�.x��cJK�9�6`�4�|6�ٕ����z�����3W�$�&��F��`��ΆG�Mtg���b,n���}�����^ƥgo�F���q��_SfL�����F��s�W�_%��g,�Tk(��لQ�.	
�c�
��:��U���f�Y-2�a�.lUK[@5� �����z��MY��9����g�N�Y�O5b�Y��N��ٙR��g���q���?�eShSs�LaV�q�Y������ƨ��ȧ�]��w����O� ~���2\�mg��냒�j�lP�z
%����L*��9Aň�%�r�E~���}��d#��q�?�m��^��Q�!��WXlxVHYEB    78d3     da0%O�N"	l��=xw���~|4c����ߜ�����]^xM���������џ�S�����t��Q�X�	�/TOA-��I(L�$!j��>�� �z�/�� 6hڏ@PW`;e�=#���{�ҁA�}�D���r�#�g����>��SXCi��YUYD����8؉t�29�0��ݿ�בks�.P#1>�g����*f�2in8��zI��9ɵS��SG�wꄩ�(��S��͹�&o
pQ�Î�w�_g|������h�R�Q7Fw��3�m�Ь�fK�Ln��0&�1d�p�t���W��X~�'����kG��R%K�zT/4��h�UB��)��CI�c{�9�;2���W��q+�/9�����l�`��L�Y�E�����^W*<�UA�>�	l`v�*b�h�B�3��X��EX]��ğ���KW{�I�y\�ޛL�d�s�"���h� ��(c�>��@9��]ĺ�����`��w�����xQ4�����庎�
����zr@�C���l-�!;p]Xw"��{���0ja5���沝��2o[R�0pݼpNӚ̙�^�hA$z���񂝁���l%��'�>�r�Y�>��o�`eq�h|���-d	���X��X� �`���ꍜp��׆�	�A��\Ԧ��>e)Q� �7])V�;�#F�X�`@�b���/�(@��.�������=r貽z��_}sIn�n��f� x�<��z�L����b�؋��!�I)�B�t�q��YR����),��P�!)���O���}��>�ҹ���_��f��D�maS���%�N����Dw�����6#ڃ�fῙ�{�pé٩@�1�73j �j)������9vv�%����q�ƈ�ƃ�:%b�;�gMɷ���8I�;]I�Eӷ��T\8�^��d�n'��=�h���\-]�}���e�}��d,��@ ��"/~���h"3�:�_�?K` $C��ȵPi6�Z#f'k1NΆ ��-d{y����Nx�h�u�\�)�Ծ�95Ģ��ЪA���3��M��
i|��~��T%�\�N��x��rj�g*��J%���)�Z�0y���.Vq	_'w�=�_t<C̢;���Ec��ي���I1��5��#Ɣ��/e��oi�?(����'b�E��5�
054k�_=7EV��6Ur�7F��C��>����ƲN~}�bjt�'�u~`f3���G���g�ۙZ4}�A�� �d�:���&�YH� :��D}Df��pbKM% �o�����y;8�č�C���o���*�\$o{�b�����L]�+��a��b��X���53�1O��Y���i��Dv��3�&���&?��Ӷc=D
����Yo�\�H�P�����9�W�Ҍrӆ�s~_a�x�e����`���������(YF-y�p*�˖���Vtp��	�A�̰�������'${W��[�g�>�07�]�̌q��<� 6�r\&2�����9��QK��K>�q5#e~�ƀ���z�H��6u6��v�E:���,��e�ar�d�au5�)��p��e	p�����|�RbY�<K�����U(Wҫt,5�.`M,�5ڄQA��-�A<��%���ļC�d�MT.�I����ͧ>J6AɌV��*�yꅋ�-w?�ׅ�Q��|���~Ԃ�w��8�b��9T�h���'(5�6�2!�)���iV��7"���V�NQn���ݠX�)��XNր��H# az��*�U�*b������C;w����O�8Iy�����!6~�(��1�a`�����"�yx�Y5\T��������P̣z����oG��)$�_����hY:�l�oT�z���Kn��p��>nS7��즏q,�M7g��U�Bt��ִmXǦ�BtȸF����+�+�ĿR;�y	�B�C��)=�<��A>���w�>/܁�ϙ��B
��`cxɜ`�F�z�}ɜ�:�qC�N�%��UpK�}G���ǿ-��5}n\�ʋ�5��b˲�6�"�dl
�����+D�b�����G+�dt*1��G9�@�V�ur݄����ٴm$����L�ڶ0.��,v�j����;�0��F��4�Rҳ:�-�O�E��y�J�֕�(�����C�g�+ �w���8��yn�'�,��Ad�W��=�����3�@F��0���S�IG#�%([����s���k�T͏��z�����&�������o������0�9�	��䆷ۮ�U��̄�5��s� /�,E8�҇!� P+Uʺ���6b�=��&��v��3ے�_���,@ew��`餥@�!�X���5���қj��������4�6�<�ܧ���]�q&�t�M[4�r�杕��!�XlFG�(aĽ��b��5c��
j�����IK����eVo�^=���i�Yi@g��F���`�y�z>�t�[��Z8��(M�Q���G�n(�i% �KAOn�Y�)�?["�{ɘ�	�\g�TJѸv���ԅ��p\�_?x�3�Ua���W�C�V���,�_�J.�����`h9�f�"�[%|�(K�M.��̞�ef��<��Daɠ�H�,"8�ѐ��/�t����(�z�����4d��y��Q��h^ ���˰�B�Z>J�?�y;B���_(���։1��:��嶜��
�v1]�k~�r	q���;.�N���[��pa1���Ij�ߦ+�J�]���P�:��ڿ�~�, 7H!��	�H��C����)��>ev�l�`�0	%�.c�S!��iw �78-!O���^ɾ���0ԸJN��^�e��O��u��5��J��G�L#:�s6
Hi��W�v�o���)�2���-�=��&\/tG�[�����&p������g��^�nA~�W/Oy�|b���,֞��ÕE�߬0(p��S�nʹ��`�+v����]���X��P�jȆ�bV8ґ>@���o�8���^��:�BŔ�;��E;�w�e���v�A_���R�.Vɨ�&�|���3y�P��~n��������@��
T����9��·¾���M��e��^Y�KnL=	`ɭ3���7ŋ�3�W
b4ȹ���rŭQ)H�]�����r%�FA8����j�7�(�g��T�źKs�w[C�<uI������`,L!���?�҂>��� z��� ;(���o���@��2�����x���zP�ͦ��bYc5i-ʜ���YL�		�o
%Q���6���w^�k�5��BV\�d!�l���5YЭn�Q����7�=
S!D�OI9���̡A��D��3�m�Ƅ���<��\d:i1�i���7H��T����,l5\�m�k�yɹ�&B���O� >Y�Z[����i�&�Aj=�x6�mL�1���q88����V��A;P!��5@��%ߙ��h��