XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���՟/��,*��q4}����u)���z�޶����s�����Pv��[��LHu'�CKџI�f.��AKY{������&z�5;��V���VV�Q�!��$ʰ�3*���4�+�»�X�}���c��������4��֥���u������՞�����2 �i�>R��%�E�^�⛳�]�c����s;�nՏ%�b��L�O�N�G�9n{�9��+������(�+ۡŽ���&W*4`�k ߋJ�#7���y�-�;���s�kb�O�h�ѐw��aZۤ�N[��xy�~a������á�x�B����rkV/CUy�膽$�r��S�'�K����a��-M�ɬ�|��!d�+��4 q̀�Z�Q���ZB�����> �M*�A#�\hy6�*kċ�B/����[ñ2)\ѯ)�����+�s�(��փ�5k���z��ہ7�����y ��"���߈� ئ�7kxæ/�v�>>�]d�f�3Ϻ~A3b8�\�hJ��z&k-Y����mG"��Ԙ�>z�%�MߑL��YǔF���/�d��w�R-F�+f����6T!,���L��;��	������Y���mJM ZA���������2��+b*̮�������&��B��'y�?�d<��Vp&@ɐ�`?��W�j˶)IT�c���-���ь���?�~
ޖ�.��"=��~�y=���c.����y��_q����'�أc���D;�C��� �Rz@��XlxVHYEB    3c92     910b��� ���� ��f��?�ިJ)~[��SB��I��Ҡ�Ԙ����a���G����Nw����Ї�5f�*�;����L�!H������o��V��c��8|K4P�N���Sqn�Pۓ
�}�>7����.U6G�w�<&}����`%�=d9�X�.)cr���A~:�����b�(E���W�:������o�v�q��M�0iw%"�Q#���F4�@�p���<�%F'ڤ~*1f/��!6os��%��D��ﮣ*eڴ��Å��'�4+W�#�G|�7G�f#:A=�9�U�!{�P��u=����DZT����\ew*2�����g�M�)��BQ��#8ɦ��n��Z�� \~�#	f�B��j�%T΂T�mu&� �@���m���H�y
w���Y��%{��|O�x!�ƧV�(]u���:	���J�k)�&��$�)�v���6���J��N�������:C`�)��	�I'�Yb��aW�-3��6w�z�UA�� �G�{������]���}ѳD�\$�o��#�ui<Z �x���M:�>�|���9S8�����p�)*�<������0O�����ŭ����9\����&p��#����C36w ���4�k?t��f R5����}�j��'kϳ�Rb��)Q�r��L4�qV�s����S��xɝ΃��f׏x&YQDob��囂�]�WS/*v�H;w�/�Y�*�H�:��h+COA\ �>u ڌ�.�ګ�}��*����Y�o��]g�F���y��>ڇ�ﵜ��nF��q���?�4��~�>e�DP���A�d�0Yt�^���I�wh���pO�r�
bӝF�]^x��HN�w�?�B}T>���2mo�'��2�n�\̴� �d�1K��2c!0>$#�-I̦ �A0ME���:���EQJ[Qi>΋�����i|��'4@;�l�:F�;� �Qj)&EB�K2\�F���N1�Nʚ~��A<�Ҫu,1xI��*�NLMD*i���~�I~�;���-"�hШ�U�>q��B��D�?4W9�K��N��ev��/2��˯�Q^"�o�DJ.����%k�`�D!Ǿ�{�?�Y��c�o�=��pzě#]�x���H�Z��C\ΤJ}�GDс�j	��>f@*,hKS�^0x������\���k㓎!���8��W��P��t�1�ɥ�"����x=wIH���)��[rrc��7RH�76Mx*�~�G ���Xtʋ�C��b��0�D�k#�j��u���]J�	~a��_��=q7SwQt��3?���m|�2Z��4�;�d���1$��������
�仩_�|@]�L�+W�!�ҹT{������UT:!hЈ�!O�ЄV��<�Q'F�JuK�ݍ�!��դ-EB&Y���i0��j1��G-�����R�s}�qod}Ac�.���������g���]��,��]ۿ��g;33�����췯*�"��ַ�<�+ �T�T*0�)�3έ\�vGO!-�q$����??�*l������c�`��qq-�+���u #L�nQ�k*s��'F
ߝi���~*�����4/�Q!�!����w(�F�U� 7�����=i܄�����Կ�p�}����4��Vܦy"�?�Ɠq�c�����dS~�%�^�N��a���h��ˉ���A4�n��|v�v�g����s�U��t����?"���4���wX��zS�8����%��܈�V =Za���g�x?��g���up�΢�-��RS�jP\�o ����'��# �wG��H���1Rj�^ �@�og^��M�aM��:�h�2��VF"���%$%#
N���"�*�#���4�m���*�#5+r��
BjE�;=���)}>�X�J���FF�F�?v�N���:z�LΘTW5�3��Z���!Ί8W˙>��{%a�<���U�(K1h/;1�M�S?��Z�F�	f2J\��V3��}StV����|נ]x�����zW ;6Ou}�LK���q{�I���������_l�V7q �@[�{8KN�w��~[QxOcM�ɉӣ"��H���0�>E
wY.��o�l�H�>R,>�ӈ^���{�i{��z�E��N�&�pN�r�?�Z��C��hp�!���/��_|��i����rS���mX��܌�7iKx*V <~}�9����pD��81L'ږrR����R�������V		�B�]����w���?�;E�e�����ރh�FWԎ�G6X��