XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��N�:����M�)���1�9� �:���ֆ^�����0"-�%�$�b��-�u6
0�2�W80ڙ���JҮ��8?��y����V[)���N&��%'�p���H?���h�5ʗSmt/�*�o}��Q�CQg�P�E��5p+rØ߷^������{&h��X�e����u�o�æ������:��N�#3�9���U3�f��������˟]�v�	]�z��V��VC�Y�h�5�'����C�M�}]*D�G�@GL;c�x�L��!�jU-�n0��4�%���d�[� �7����+����ַC���絑e��O���65:��a����Fz��]�WW=c��$������I|x��r��=�ܠ��N<v^�����+	�!o��K�2�_I�����L�{�U#�<���X�E%I�H��GK]%QB�\L��A��la�e���1Cć�����Yڴo���q�@�v8��!��o9��X�t�A�����to��zd;7QeT;�>�)ca��i�^�Q���azY4� Mx��X���U_yWC?C�Y��jI ?X���A�
v�u����?��;m��T��=�#��8��f�b��~D�:cs�~��-��2CV՗e@oy�4�w8x�v#��a;�*):��0/S�|@��SA~�,@���M}��մ�3dW����/'�ZД����a��z��ۼ0�3f�&���E3аT؈�(���,,/�:\��}��z��.K�^=������g���8��/I"XlxVHYEB    2816     5e0lw���,�c;���챛CI�Omq �XJ�ũl
�^/>�����am��;R߶���Q�\O����E�ۙNЮ^���aD'��x Y�(�J�+b�(�c���M�M5;䙏p������� x޼ӌ;o��0K�/g�@��`�ҷ����[�~�q�#���1��$�[p�YK�4����p���MR���|ۨ��n��Z��O,��r�mjFJ�3sE�����͏�x�F�s�4�|�_~Ė�Qo�{��]V��G��BeeJ]Y�2aeH�ǆ�Wvbw�#��I�3R�O�������NEr�b�C������Q�!�k�]�X���csf���*j#!:���r��S��p���ѫ@
��c��Q�h,Dd.v�)No-@U��"��r�jK��v<�o�5���|#����� ���\j�cg�\x����Fg*�g/��2��B!!�� �0D���D�o2�6�G���׻4��9�����9$f��������m�#xp�2I�Pa5Q駠ln���qȖ�9��K;�o`��H.�;);Z��jġ�o:�,=?7D��_a��Y�ʇ�yZ�9X�S&��@{��ho�m����^|���������j��Y�ڔ����G}a��9����_1�
��W�|��^���8�2$�_%�����[/��r ����^����n��W��?��$S�`�y$��}#�{yMZ��c[`�F.���M�i�N��
h8л�U�1�Vb^�)I�ti����:���@T�=�t�v,#� �[��y�;�4�c������X����@��a��YK���7�4��Z|ْ:joٲ+��� �,�}��l����@l�[P�Jbq���w)zH�t���񝌈+U��}X c/�?8�O��|N�c�@fII�;�Y�P�jp��,��F�⋗'E���6
��g^n�潘�45���~e& �]���0�]]FX��U�dG��J��=�pפ�/��x���yx��Ǭ�e�� ����l,E�rs@+{�:�p�і] ���>F!'�}̷��I��N��?��R�ͲQu�F�t1揞<�
r�iq/����ɕ�\��Лn�_<M��Y�d��+8��$n<���3�����J�߭�w�[�k尭� /U�1��p�^��6��W�{�$�aAʨX�(��a�e���;hY��4��>U*��7k2Q�N�q��V�R��!���m1��`���#�&CF�"R���_�x��-��k����x�s�mώmf�9��܀�o���*���QU�]���3����꺿=���b��H^���ކL/Y7m:�`S�K-�G���#��J|=�qH�\O��0x
�k�q�w��9��؟$J�B-���؆�������J�	:�V�,�N8@��Ȣ��Ak�,�S���"	_�.7D����x��ؖ��;����M\DXܚ\<