XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���s�q摝F��xXw�l|�.�3����YG�L���ȏBN�`"�D�߅ǀ6|jps��}�i��X��]Y�@b�� Vb���EU.�昻T~��6�Vi4��7��x�k�r�y�O����J�Mqv��"
�Ra��g�\��t����ɨr|C�}�"��о5��gy��������"���?��S�nMe�nR?����ג��yn�-Ĵ�11�o<xғ\�<��'�a�EM�^��Y��]<��OTl&��)
:�O�l����>�gbY���>��T#�y�����(,�{�O���O��[C���'S�ǉz���3V/ݐQ1�lY��
�70 ]�#�� �UD�mObL�;0�vh�-1�=�Z2���t�f�mas�Gc����/n�����$AT�b��U�p}��*�?m�|�1�p
�Q@�c����e�0b��7l��s��[�Β; �C�6�c����͋�R��?�lvo(OM�������7N��C�Yd�ڝ��=��K�=��Gd���/�wkE��&e���f1!rV2��3� �XM���*9��ü"����d�8����CF!����˓��eȸ-�
E�����u
��\�x�\�y	�;;��K�.�HG��������rWJ�!C�w<)��ă��K��;M8
�X����I�?��/�4$���������Nmr?���@�M��nI�����'���L�靿^���xd˒2�p-���S~D��d�#]l�g��2��GXlxVHYEB    156b     590�6�K�e��Ri�������D�턼$I�x���ƾ�u��"ZI�w[�܂,Η&���������P������[��P��6�mA�]���aȦ���Zs��W����Z����HnA�/d�Q[�?�A��b���]ﾌ,>��-�����X�,��Y��mv���R>������ͲI��L�_֔$>��t�����aw�bT8<Ț�/��;7���Aщ��5@ڐmh��-N��MRo�-޸����0 �ʼc�O�WG�a��v/H�f��?KF�w����g�` %�L8ƿ'${Э�S���tUY�Fh�У�D���ͻv�u�ܱ��߳��m� �I�6lV�L��Μ3���8�@n���V�KD[B��y�|`�~;�g�H��9��1��	k>�u��j���wT���J�����\��s
�J�u����e�f�!�yX�EP���w�GsQ,z%����[�:��;)�s��uD%��Վ��s�}cy|Ò�g��vi�F�Y��g;��c�k߻��k'�F]��%nb��SB6��9n�#?I?F��Ǯ�(oL�=b�W���82�W:�R �;zh�S8s�t߭J�B�Jrx~}�#D	��IG���\��F�~�nV������Z��� `>�NOˈ9��׈�L���&��Bpb	���*�Ft���Á�cZ�"FJ���/���k�*8��x�RÜ\&=�?��"ֵղ&��*86~�~l��@��v�a/b�~�7�2g����[n��'���p��-E5l?���_��ǀ��r=�?֛�G� �?���wc��_��N23X�
��#'ާ@���R·)��+�[8��n]	n�=/d��|
e����`���wp4>��(<��%�Y�P��&*�0Y/<-p>v��gjg��Q�wqr:��5k*�)�I�h�u*�@���*4�m����p!A�mo�;j���B���gl��D�Ͳq�[� �@���w�����W���(��0谪�ב�^9�(4b>/�1"T���������$h�{�[��6K'ea�상������vS��(�#>����92�Ό�r�XV��E�k� ��:����{��J�4��Y& n"����~Q4�ͮ��ˌ2�"�2��w�`ϰ����٢&X*�-���0e��׻m�$+r�/)�ڜ#[�8���ٗ@�f�Y�s��!��ai���cm9w֌�NGF�Iv+���@Pǰ�&.8��q&gsLI�cR�6��R�QT���\~7j�s��+.W��F�r�H��]N�6:'>�*�Ñ��2�c �G��g�Α�9���[�_�M9g�����m����E�csF�RU�?e��F&����7�P��It&l��$0^���94������A��A�ع�;��f������