XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���c�OŰ��[/�a�{�������i��<�(��6�߁�O�M�l�!����v>�¨
U!i����l'׽7p��������'���I�^���b���9�Ӯn/Dkft�>RR�~`.M���J�z�]�#s�i8���o�"t��� >7j7:rdr-J���8������p�KaSżl�c���.�f���������Y�g����2B�z���~Y=�������~Ya���Z���z�%��V>�o.��RJ�9F����\�{q$��; �X0���o���/YE�:�o�ւ勎U��.�G}�T,n���\h����S;p���e��a�3�f�p�ܢ��2;~��*�"��V��;qpMXlHV�����I��M ]o?.Q�f�+�*����9/S�t�iK2x�VT'�6�Ͼ�c3�w|��X?�hA[�S̑O5	d�է���i��|{0���wUr����)��
ڸ��)��w<�e�t�'�H���[%�Nn�gٰ@KSĬ̝R�9����Nk� w�Q>�����>e泼��9�����
Cڬ*Г�y]��7L��#f�^�z�"�t���뮞i�V�%�+m���&`�F¾CӞ�Kpݎ�����b(4�%���$r���0OO��]a��W���U,����%I��Q�/�;t�RI��Wt�Y h����A��Y+���Ǵ�E(�m���, z�l�PGÎ'�9(�~I��� ���[�/�D��2��	��ܴ�ZXlxVHYEB    216e     8e0C;���:����#yv��ѵ���<:�� ���f��I��kƷx��T\�gN�ſq�>�3dzxm`��+Z(��Y��{���˯��O���`q��%�h����h��J��zN�]z�1F�"kų�R�4�˩�V`���|^�	[e��L�cAf��C�=� .��+�M�hZW��-o��M���L�Q[|_�wfF��lm1�@A���f��"]!��Hl ��d���1�6R\u{���Z�?Ѓ��P��K�!�C��Ńm9�g �^C�߾[c�eI=������J�k�˩F�T�7=VN�W�[�qb�f@& ���S�L��Y�2���!W�8�`:�}j��1��p�ی�rRזuY��5'y�ʜ&3S?5����"�py�Wɏ�������^JS�_�[I������֠ۘ@�ش�������	\ V��v����HY�Y
B��X�J�&1��(j~�0G&h<��f���H��1z\������O8����$��6I+Z��,���MYR��n��XBZ����Iþ�iq��K���/�?چ�����Y�*��LG���)Ɇ�ܶ^�L�ռ:ё$U�`��y6�J@7q�� Fb�g�U���+���|�5Ȱ���ǽ�e,�ϵ�]\���:E��R}�&��hiM�L&��G���-�(�*��폙#�n����̡� ��_���Ɣ?��Q�"�]��-^*u�_�s�+��0gX �.2�AYs'7�ݻ��{k�5�����n��8�~��m[(�u�kBM�8������ʶ"��5�b�8���ec�Rp�k����d0�8�ߧ׈@��|6$���#lx��A��^.�=ՐΥ%�I�Ν:�K�Dq��Za�0�� �*ƕ`�Z����7�����_�Xy�Z�l2^��M���&�K¹�"��l1�?�2Y<�e?Q����Y $,�.Ul�/�)=Hn��Z����L����̀=&=��Q��@#��q��nG�f?�8%x�O[�;Gd�Y���^Y�ׅ��m��<�df%"3��M)�`��\��6���3�uWd���t^�ŧ�0�Be��d*�R�>�d�� �e�Nh�6���	�@R�@�F���K?��=�^��oI�6h�A�!چ`���%fkg�r�e7���!��8af��$���32���Q�RA��j��6W9�<��_�%����ʫyd_������k�k�~�5ÈX���
�s͵�zgR�¬����Z?�2��E��
6���'V�QT�ly�xʪ!����h����]���!&�IMd*����ff��M��~�`��ɤք�VpBq�{��d�Q3��۳"G�N�B�&؈��	���i_��PS=J@Z�)���T��#p�~��##���B�$�^�ל�v}�l��'�ޏ��'p�ow����lx6��ޜ_ϞN��^�+�%�'��qK�MF���)ȴJ&����o̮~���`��P;�󐮮���2�%ht��F�_m�l8?��BBy Ѧ3�*��GKw��9�3TK�\���\�_�U�):@U�>E7/�+ߜ>�0����ݑ����R���\-�$�%V�M� ��ak����e�f�mUP�B�(q�d+�i/P���£�m<�N����5�ձ�B�Gπ$X=-��)[
پ!Q�}��*����SUn��:�H�b�!0t�2G�&& ,U�*�� |h�o�%"���➣��O�Ć���Mw���$% ��VK��N�TN̋��V�Z�S����06)�e?;�d��I ��Dh0�p�����h��B\8��bj��Y��4vm����^\8/+ ��!.<1m�C�B���ة�[�,e/�mGT0��
��om�SCi~r��2ۺ��l��qy|�"�̙�5���4�L����\����F����y7��p̍r�b!�����4I)q�Vs�d�V��Xy�O�P��z�+�o�^�"BjkT_s~5��A�	V�5�B��ƥ��&�����g���|�|��g��I�bV(�
 Zp|��u��	>��p|<`&>��:ns�"i��O>�em�N�`�pMM� �+%j�-ŭk��$f+S!���f��0��͊�Qw.ƭK�W<	 ݨ�~B�^ʥ�Xo4�#�}ȡ�8�]>�P�+`��Zj�&��y�еd�yr�g���hx���	�-�уf�[$�.�}L�1Z+7�