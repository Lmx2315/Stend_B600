XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��i�U�����P��Q)�,~�U.�)˳@�\.c"LU>'P8�ɝ�40����W'~)��V~��i��V<4�� ���R=/��X��,�T˸���_�b������Ҽ�Ac��\��y��I�yl�/�A�vv��C��@��]^[�!ƽ���'ӽ��������ߦ�����Ưs`b�W�O�G]���ߗ'�ߛ���:��m���)�ey�RS�ǖ*�O�\��b�)=��_V_H��'R�c-��<�Y����6?�ٜ�����Ϡ41�4m;��{�u&�E�gp��qs��H�E����:�`��h|L����K��Y|0��#R�Y92�5k{H���EZ>��@���o� L��+�[���� џU��3��R$f>��y�)��Do�%4����aj��t�	�^�ـ<�I�� ;U��E_�5�Sq'n[��g���.֗A�87�G
��DX�_����C��Q\�VK���1��ϥ��%rPV]���;E�c�Kv�a+~Dh'r[�{�����)@Z���Q�,���A�)��"�z���ܢ���(��(���+�2"��M��������SE��$�X�rE����:C��1[𬏞.��R�gZ��j_�tF;�י��O��ֵ��X�����rE�� �S�2�/PT�����o��5�����2��U�iГs��*������>F�}��[�#���Ǜmՙ�GA��@�Cq<i�@��e��Ү�;O�đ��XlxVHYEB    fa00    1390�r���XU��dL��}(���^*{�4�eK�)A��1po������Y�*/�l.2.���V�9-��.4ō��f���I2��5�qh5hZx���1?�w�𪚩�Jj���?�cxD��b#�pHT�~�Z��,����3DP���N7i�Ҟ�~����'���\Q�&o��v�׵
4_�0�����i����˅��GT�7:"���㦲o�����E�0���o����:~WQs��y5��NSH�L}�0Î�/�+��]s�N���:PS��Ab�TA���1�u���ԯ���O!��~��/�u���c#؊�{;��cBؔ@ڌ����
�ǚ�`z��=f���B!�;�H	.!F	�칀��.Qa��L��{?f�G�~Nm��A�%5Y!��+���ʢD���n$ڃ�B�B~���g=ʼ:r���5�M���V��jH�S��Lc:M�jU(͟F\,��V�`r�B_^�ԭ�	v�	��ݽ���(��'d�*K^y,�ЎG�Y�}}\Ԫ�f�7eC��0����a����֤�E^�&�&)�Q�]+���tj��e��!rP`����Kz��[��RV����5���{}�֮�����P���S�����]���fU��w��ɻ<S��_J�A����$��ni3А��;j貉18d����9���5�_�E�A(]TԿ��!&��Ћ9��"8 q��ѷ�x�\�2��ߝ�`{A[��kMĬ��I�t�[c�rs��s���K>+sG!�@X��F��ժ���+�R��̿d0
����H2Ez�|@U��^d�
��B�67�#	��M��+6Pq ~���#k�M��#�s�7=,��˷�4ض���^��b�4T�g9����M6J�j�Ho�B�������|\r3�R�w߼�Gxpv#܈S�4,�2��}��!��=��|Zt
��*��/��lV?��ݿE�.T�������=#V�߄*�������T�(��A����z��Rl|$Y��w�Tei~�O?-Z�D;� 8?�ee���Wh1S�d�~�Z��.le�r�uA��t����:%��J�F6-�H���2� �_�Oi�ށ(	
UwטM�  �f)�q�˗*Qq�ǵ��#��C�T��g#�G�Î[v j��)�����x�4�P&ނo�k��s�Gϔ�\��,۹�=��ǃ�x�� �ї�N~SG2ӫE�R�T��3�!�����ܫp�6��s����A�W��k�i�'��W��r5��yS�7�W���7}�����<�G��INs�Jư�֕g.[a�I��T��n�z|P���+�;�N8%�U�9��I����J(�K�0'����[)N�F�[G�u��Yw�(v[�&� ��<�=�/�Ϳ��萉������\�=v���w��x1q�
���63������H�R���~O�d�+ ��B$�e!:V��O+��?��6D[�!������K�!Ňc�_�H����(���/�=��C�:��`��uL�����k��V�8������d�e�aO$���4�� p�F�׈�dEY�.>��K��x-v[�<�q�Z����+�e�\i��{���)�3��?���&�*�U�X$.��Y�$�ݢ~����(W?��ڔi"ɽ���ñ�i��CW\Н�p�k��H���yU�<�JVBo�
@C��P�ĕ�a��ATD�1�GuQ�-�A�-�RW�����;fu��s��i������V�!�-Z$�=Y1¦N���j*/7Շ_�V�jĕR�/ܾ�Gh &�8������j�	����W�[m�aZ^@s�+;/c�}¢�|�"֡h2����-K�E$!��euF,�z���k9 f��j�99��:N\S;H����RI�<�^�����^�"kˀ���̞� [̬��/r�)��'I��QW�߁��
�$���"��9���(��� ���<�'^��j) ��x�N����Uݏ��G�3�erQ0�I�Q�i{�NZz�d��H�m@�UI� �O��~;x�;Vr'����r�ۈT�1/���gy阊����X��%9f�[�E���j�{r ���Ԍ�/`�Ok�}e�k����5d�-�q��O�乮��l7pA�J6��XN��i�-w���z&�~��
�#0ꪒx��3��+����_�J��[�ʬ?�j!Z�x~��o� ˂�h�z����֟�iJqE���uqAEϤ��`�G��Vs��I���ܪ���ߛn[�j9�y �t��x��ib.��Acd�}�+�ICHo��2�[ح�Ty�}�����E�x$i�y�
w�r��;��#�}�9��n���ָa�-:�~�9�'����B�`�\ف�/%�c�& b<�&�<:�2�k�2#/Ȟ�1QQ��	Á5���cS	0٥8$k$2�Y.��ߣ-a��vf��n�*9��bh+"qN�B�*� Hy��r'ԉ��d��{7�3,��h��7�?}�_�	_'i�O�A|�תG�N䚴�@�C�lw<�����j�<�FJ�qI�;l
`�Ս��~rs���L/8��������X�g��֤`k�C��-���^�H�8�X�3<�4�xQ��[!�J>,�d��E�����N$fs(�0��h��h����:�{�]A��k��ɯl���$�5�(]3O����q��H�T�� t��!@S�U��=��9N�RY6��>~n�����O}�|)�'l$ͧk�ECP�>0���bằi��6m��}�8��Q���C#�ďJ�]����
����(�cU��X���	۾
��/�#J�����V�B��oV���N*Y	3�����iۦ
&h���g�KF�����i�B�I�홃�/�̔�xP5��sW�>����:dM���Y�Z��B��}3y�4�Al��D,#i`�gg��A�]��$
�Q�/O�k�H���p"8�7$g�f �I�?�p��f.�O
 M���T�Z.X��ߣe�Wa+_P%��EV"j+η��/�G#a���#���!M�W��2.t�s/��2�ّf���7��q�=��kTUR\6/*/czY�^�3w�y����*� rM3�0l��E�%,�F�y�!,i���#�u��)Fy?[���$�H%�Q��C���O<�Z�u3]K.����4!��ss۲�����o0��+�/�k�%,���eQ�J-\n�c+K�8e����1+�FV�Ǯ�vKQ��X|@dm�u��R	���
����2��(c�5�^C��B��Mh�3�1-�9[L5�~���g��?�6��Ő����>�%y;�[��@�GQ�.K
$���U�o1���U�7�_��uQ��B-E�����͙����3�0jj�V�t�"�Uo��\Y"��/ކ��T��D�k͒ʙ"T˺���2�0Af�� tN���*���� O9�*���mu��P���E%�s�0�;O`yn 0̡�������\�8���G@%H��6c�ļ{V0Z��f_+�z�܏j�
/Enf�;S	7�d1�X[.���I�-���j�6�6'"���S��sR�{�)]"����{0��-t �C��w�)�G�A!vd��Vڥ!�l»W5�I�`����
̧��ȄSWĺ�H��{� i�./lC����f����$���y���@�s�k��9r{��wJ���}��wl~n-|qH�ȪD�}�-��v�����}�Q�#�!�l��A���E5��zH(+�_:�շ�m�➶��[���	9��$�sM�%`u*�r}d������+�}�ԋs7��d�v �v<���X�ro�p��;�����H]Xj�C )�� -��8�Pۍ��yi�4����������i��z��;{�����a�T9~?�B���3]e*�J!��Ե� D���� H`�r7p�6��KA��ie���(����3u���a�.�yZV��7�@�f���9�ڌ���!�r�7E3���v~��'�����?(}�v-ҁ�d�!��ۘ��R��5h���A��M��C��8���f�YLL��lz�jC�Z�Y�׃bڵ�,˗�K�A	���	�/>�c*�/Oi��D����tE��v�S�%%�,�s7�d@A�ƾ
�Z��=u~��wx�L�i�3gX��Bx���[3���S;���x/���0�:����!�O�s�W���{�rr��)�
P���]�����=��K4�Rvǵ|��	�hߴ|�K1�|�"PKp�C~���6_� �@j󈞖u�]�y�VE���ڐxF�|��a�$�O��]��a!����u��(م=�S[���'p��7��g����Z&$���K��5�M���ߕ!B�Av����.ڮ����g�>��@Psb��P�EMOFh��N��c��U���Ǹk�X�Kv;S�h�š�u�����ܤ�����5a�ה.������`i��5�o�ȸin�DpMK��dT�.7b�{�����Q�ϯ��.*����v�5SdJ�R��}�+B\��m-� ��c�J�|.J��F)��\D�#�˝�ȁ�*,��]��@��2����4.~�ծ����҈����	�3-��q��1�eC�Q��E��r@׬�g��8�Ѻ��俁g�����[7�����awnB������jb�6&�߉Ƚ4P��#��a�"1����|{���)BR~�|ƥ����Юn�wC�zu�b����0��8n��<ʹ��゘S�}�3�#/�?i4��wL7k{�����yM7�ƌ�K�,��D �/�!$��D�2���hU��i�[��C�gW�Pݮà��R�K~'q-�<z�It����RP�qJ���R/?�I�aĶ���jl�@��~�{)L��~�A�.x�%���r)XlxVHYEB    1193     3e0��]P����{i=.���K�k����#I�'5M۞�tLwW������Wup��i+�I�{.�&t���7&9�
=���w��;��ާ?����EΪ���d(�uv$�5�ھϨ!��9>��|�d꼷Z�y�OL㷽�k�!Gz�mk�^����.OO54ZZ�}V_%0��!�����������s�/e�BV����/'�\|���/��b��|�w/0)�S!%��>{|eQm�>X���ap<��y �tK�:�eD#zq>5�����]�1�����2s���ƎR�h�h�5��[�"������_�G[��Z��P~ވa�Ǖ<�R�e���Jȯ�L�90H^#̱K��H�b�d(qC�%�XJ}�l.�US�Ŏ�k��ZJ���5���U��\X�fٕCg���<7lcV�|���Czrs4B)��(����U�-��-ϊ�QS����l�V�o.�C3֋qV7T%�Tkk�1�f��СS��N兑mP��FU����/�׎ׁ���w?�$��N���HM���E�)�a�_���i|�P��r�[`��Zu��ʹ��A����(<�R?��=��o�og�09�lȳ�mx.9SD�aX4K{�r��^�Ã����:M�D�Z>�MJ�M8?�ʀ��ʨ����$��?��8������u��x?fڟv�LT�uz��ĭm� X�$-f�1�UĐ�K%|��Q8ߺ���2�����BFP'V�Hm4�����Z|�: ���t$��_	Zqq��E�̙�}B7��z�[c�uRF�����R�2x��aX���-R��܅HP�AH�I����P���n�p�v�y�0��)�`n�h�m�9_w�Cњ� �,t����C���!Uѡ~�Z�����E&�S���{T��Q�֕�W�����}��(8�zT*�U�k�h��eR�����?�I���T^�v�>� ��%j��wK�+��6��_�����D�*���Bu:p�w�