XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� � �SA=��1�K�(z=0~��J�A�@`�l~������F$�r��֢?GWك�w=���p9�(�~?@Y&����$N?��cpXG(��	>��D�z�-��,C$.���Ȱ��/Ad���IbL�3r�"L�y�Ŝ<Ly2��(��"�dA��j,D�������s�`_�;���W�ېQW�Q@�k����I>��[ȋ���ϣ�j�p�4�����u�ClL�j�K�_V�ȘTh� v@'�5��sM�2��ء��S)l��M�?w~P����fI�v��0J���8�/�/�8�(5O���/��|AݠHq����`���4����h��B�3f���ƴd�e ~����f����	TDC4)��K���f��@p�e1�5�~W�<y+%s�T�4x�j1 ������6h��#=F�ԀQ򃈼���8<��<x�Mf6��<�_���@9��Z0�5~�f�uň�5�����y��#�蠌�C1P�� g���\�tg��-�[S�s�H:P�]!�b?�{�!�pE���3�3�B9|���9����s�]�@p������=���k���n�?z鵑����3Km�:�[��J
U5�5aA���~�p���C�n@��TS�*���VN.?5�z�q�����1�Z�;���d���[FE݄�?]�~I|ANT�����fT�0B�st+�@}�4���iɣ��G%U��I�<�pu�6K�7S%�}KӔl�}��5XlxVHYEB    1621     410����*���`�fYa�W��&�@$i�����6�*�f!O
���~�GT���Bh�_��h��݀ϝ�+sr~��Z{Kݼ�:���Ƽb�\W��Ϗ zU9@���Y(�׆&�����Nx1���#Y�\��~�s��.4���0Ka�v��:j��2���QkՓ�Bq��*d�'� 
֘X&k~���l��@�%�^|N��4y�^	|L�␥�����G�]��CM�m�O����Y<�Q,�B��+)�k�e�0��T�v�� �Xeg���#`g��٫A�Oq�o���B����P��ӿA_8��m���@d�f���ϵǥx[5�ak�Ğ��5\�LAv� �Tx��@�д�+�����L�n%ء*���>B�t��թ���ƨ*�\K����l�;�{��J9^��!5��PN.�='�.��~|����WM�5�����/��b��s.�� -ٜ��zZm7<w6��-�+��~����	�R%#�i^yZ,�$��ag
G$��T?�tF)��2�
�[�YTtx�-2]����l/E�+eڸ��T8�<���dQ1΀|@�o&��U��a�q�ڠ�-+-/�
����b=0�&�#3!�x�.$�CJ=�Bh���,�H���I̎xĻ�%+��cc���C�jwΖ�E���5��O+�܋�~�pg�O� ��`m#�o�^��!'�#�����.��H�Z�X=ߖ��Ԣ�ޔ���z$̸�f��H����W��&Ig����X����D.�4��7���X�=�(�����/��q���JG���G��ƸuV�i=�f���u`3���:�c�T�a�8�T�<�8��S���e�/��K��8��sބ���M�\:��Q��<O����0�}�b��6i\�X5io����VٮH@<7��`�ׂ�/����9A��P��?=sv9��ܟ�qm���Г3�r��NAw�z�A*�.�S���L�G !�v�n�����m3���x�L�Hќ-Z�e]c,q�ˋ�"���C�@ն+�l�c=���