XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��kx�A����9�@N��/#(���t^���p̝�/)��8!G��8���5��^~[�I�0����߃Mf��ث��jz�c��'�Hn։�+H5.�v׏~����%q2�D'
`A~�m޽&�J\�Hc*��\�S.-�'qɒ�fP�\O���(�����ݜB��0��/2��>]��w�>��s��@Ύě��������>`�߯jOC3�������|2�bX�!�_��)W@���n)��G���}$ClA���������qf4�t��|�C\j�0��u�& /%	G]wڝ���a�n�c�P�M���#��g^�1(���4u���^���"���|)���G��zh���w�����b���}=���5�<� ���d�	2���ᕨ �A���� $�I�J8  E�%u;�-߳���ڞ��R+��}V����fE��W��h�]���� _��鵂ߝ���l�	_� ��/�H� ������Dm�(��Il��r�=�~�*M#�[8�8 ���3~B�=!�[Vwi���s��2���83�>lT��DX�i�I�C=����,a���#�9��tZp@q�Ú��r�`٥L[F)�|R��d�ϊ$&;�Pv�5����XHl|�+�bq�뱂���z���c)�mˬ�
B�8�h�j!ĉ#�KI�͓�g��V�z��h��I�c��#���X�J��Ǒ��:��RS^N���	Q���~͋���	�E� N���3�������^\XlxVHYEB    1ee7     570�"yN�	QV��X{s�L��(�V7��Q�?+��C_}�ĩ�z�@��	m�'ީ������
i�8-��3��m�ؼ�S~3�:S�q�`1�V���$��UDc"�E|�Oy�[&!�z�nx>�<��������S��^��`,��=�4�����_���5FAeK!`���M�GB�\�k����"H�����}Ʒ*/!g�w����rjMR0,c�W:�_&Q�O\o�_�LϴT�"9�g^�nھ6B�K}ׅ�����6�vb�p��K\Ԧ�Z��2�@wK�;����I
��C���@���1��ٓ=H���}B��N�^�G|g�g��/U� c�����8S�J�'1L�̆l�ʤ�j!'>h��,�N��m���x��ZH�\ו':�[�uh��{�Y��@�/0�t����×(��(�~mE�n�|�Mtm��,����E���/ ���ڏ r��Z$��
�lo	�z�l8$��Qv�� Ӝ�5��.�+URDt!C3-�˗lqyo"�S�8g@�;���~���pGeik�
!oJ��4�ǖU�
�\e��cAKa��2Λ��_i��b1�pD�	��F�� f�Ya���}��G���<أ����̷�]�P��୳��PX39��]Y����NPG 镑'fk����g*��L64�ߺm�	i�P�[M�0�&�5���q��`/�q �ys2�{�\���5|�ުԉ��yL/��jB��1 ���Ac��ƈT���#n��Y3{ѫF��n�Ox�V�w�/�=�%���4z�q�1O��]OZ[�ե:���s�X�^��>T=�ɠo�(x�:��C��f��!6R*tg�Wi����F�P5ո��Q���Q1�u�,�*�5��a����A�L�ßl��R����Cu�#� ��J�]��g��;8GQ��v�֨
˄^�Ã���w���ӣ�z���WvjϷG8�&N�)N��r�gF85
ϣ��2�<VrtQȓ��8�$}�/؁�JfxP�|4:lR	�+��I9�,�	�R�wƄ�@����V�~z�1�h����{W�#ʃ4S� }��K�;���$s�N��]�e�7%Y��.���Q�-�䗅�����2M��D�����-?�:�)��&]_�x����SA�E�!D�`�"�*L�S���#݆v�e!��'].
3i["���]g�d;�ubƲ�#"w�`�@r<��\�Zx1�q!��1{��}G7�E��9�2�D�ٌ]*�W�C)��4�.�	hb���rw�b=	�?0g�6�e۫���2mB`�s�0H��Њr����'��-�C5�L�E_*UY����,b�sNp�#J[��