XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���7�f0����dJ
�l!�{���?}���!�V���0%dih��w2L�Ni�P@�ڟ�.�g�<�E$�b�83-H�|����ؖC�������d���epw��"`��B����1\A�D8�p����-�q��U�n�S� �9�{���?�rB�C5(�JOO/�\�-�Tx��bQ�N
c�9��Vs��b�*��i�V�YF��T	kT�_�ĵ��¤��=��[6�:\�kgĘɛ�4�|�@\2h�h�y�Jס�.[�dä �g��v��Z�!����cC�#������ ����V��i���!�C�#�/�����#.�F^�	P������5ΜTh��5��w��vR�4�5	235��-��W[C%CyS���/^2�*:�2����5�q@�N���u�l���g��#<X�#�_���u��Z��I��1E�;�_����Md���Ի��jn9�w�Ε�X�b9j-E�X����ʐ>m1�\5NS���k�-��}_�$�C��ĉ���kib";V�Y�$6�ZWuVHwZ0G�i
��ۄ�.{z�C�g�Ԧ�f��ӛj;\�1ͼ����Cl?��|�bad�B�OeX�ʻ�}Y�$�������p輇�Qq7�β݌��j`!b7�ƂݲL���E@5�BH��\���4�#9:���ZM�,/K������Ē���|-��n��KH���'m�|�~9"�(�TK><�(3����QϡJcD�T�?��,'���%���jw���v��XL��XlxVHYEB    5ff1    1040J�������g3X��Q����[��p&-��	������|��1�jt�^F��	z�)6I��&�2���d����,�֟4 wV3K �V�ٖ#����<��O��S[xO��l��*�<&��S)Xऐ$Qڸ�7���ȱ7�̨����IC��Sz.7���F�ċ��6:ru���|!Z&kpu=��v? ܱ��p�| �r�oC�W"�\�M�!\RۊѺ&�l�����V_�Il�P�Pe]�>)�s���A`Ќ�@�k\���'3��z����m/�ؒ�y�}�0����t�7��P Q�~�"�%7y5s��K���F�W�����`j�!����w��l2�و
�7�cN�\[��D����ō�g�*}/��^/K�N]u�a��� �&���Z�D�������P�Rwj�B(lZ]w�F�������	� ��}���^>aSl��-j��ӶH�`�4M�t[J���4e���N�7]A�����La�����g	b��P�!;���(y��i�ޭ��ٱ�HuVM�?T��5��
������:p������wZ����l~*�a����H���T��n���q�?�A2���NӬw�<��W���2Fu��$�Iw�WT�."5�J�b� �6)n#�)�@$9�?r;��A�D"�e]�Y��h�y���D]�F�D#�s�8�R�(�[�Ҟ�7����=B�OR�'�J��I��9y�h7��q`w����NqWA�U���^M��2;�e��4ʐE=�����d�9��Ǧ��m�5�K��^�3�,�/υ�p��]�ܤ�qb7���&C}[8?��xߍ�W�\.����BYJ6�K�����sr����Q�A!�����<#��d�:�U�]�6g��K5��U�S �z��}��J&/����E�~㞾��fYQ��9$iC�!�*�*,{���ڒ�T-`�-�H;P���nx ��?YTQ��.M�i�sb~|���l<��0>q}�&������(�^5���Ń�}���X�肧�>J!�Ծ����[�� J�p�i�ԕ�I7�Y������A�@�"�M�%d��eJ�\bgn�1V�NƱ���2�?nق����d6�S꺓���栫���U�#�~D��}U�)�N�%� %�Z���	�j)�S S��¯�S]������jѸ���Ii����@�eo��7]�mbǉ�4�`'�3�Y��Z��Ӓ6$�ν�ȧ욤��&��{�r�R���yهZ&����7Z�Eh�Țh�u�
uN�̫9�d4Aa���<�OA�b|��п*GxGL �,:>P��}p��el(G�]Sµ��1�ㅳ�u��F�$
�f�j�lL���2}p�ma�UƛT�o'� (���؞8�A��0݌x�J�J���c�/�+��Ùh�_q:�(�宅�T���zu�v���wsmXܲ�MO��f���sD��x�����T����e�r�h��p�A$��B5�гә�nV�m�5V'�6�c�}w�U/���Fr�>�51Pp���QFD�V�Qڄ�U��] ��2��A'���H���vעH��J�q��m����7	m0��|m��j�|N�l^�{{�LR�oʸ=�4!!U��mH7�4��Np���}gR
������F���9g���*�o_�Po+/�|�i~e��:��հ��rU���2ܨ�q�z9�Zh	!��˓�yX@�I�x�/c�1;$(æ����T2��+3�}جZ��'w�Ü�ӥ���tZɍ����f�e�M&�:T�O���ᴊ/��_�.����B�zt����4��:������'�k2�)��F�e�"���<9)���zA&�/�L�4~��a+���"N?o�+��J0�܃R�O�kR�SK��(�i\��;�1�o�˜2�G�q�2=������ ��r���O��K���4ލ<�@�@<7$V���5�ꤡ_;��Y&/w�v�z��Ճ>sBo���|a���.噙�W���,�m�_��N
�vE�7����WѨ8Y��������9� p�#�&Z�_�QrxI:�I�X����������9��,I�Џq��V>{���گ���s>|����'x��2}�T��Dؑ �8yx�7�U,@���F�"I:!z�0�F�}�'��Ii%mA�Ʈs�a+)%Vc�d��O���.J����R��>�\b������¡4�q������yh%/T�A�o+��)�Y��s�q���v�n��D(%|�0��>+��%��ض��U��:�P�88l�[%Hu@4g��V���*�����*]~{�W�Z�PkYf�L�k����S��#t���W��=?n�e(rt�����V���I:w$o�����WB�~#�ǈ�೹����K3yC����p���^�ֶy��[��� O�����9�o��PЂU�_�t�n�<��Qŋ�'V�ίl�6SuN1�������I��r�_i�A�Z��qc�V��b5IT�f�txT"�	/�g��!�!S��K)3<�-���J��|�L��xTI*�����Y�88x�vl�O���/��dĉ繹�|�^0�3�~�W�e�HSck� �vPLJ�E����!��k��6���݁���������jy�A�>S�$yޥ�@�n���{�~�W��������|�B�8�U8݇��w۽S?��������VR^P��� i)���s�@u��.L�� �V�T�"�jPB]���6 |��*�����	r���8��'��O��R��D�3�	�N:�-�y�'�����J����/���_��c����Q�8�/��P6uU�]��G���n�d�����Lz#Z6b����Oy�k-�D��)��Q*|�x���T#R��/PˌA-���:��6"�>�OZ8�;�>���v���ލڛ2D�<j�6.n�h֋$u���t�?��n�*;S\�9bV_\�����N��eds���g,yO���T��Q`�&y�#P'����\.g�\�>��|�����𬲐Q�k�7]�C#��������S�����FI@i�F��E0�g��DKi�$`�6���^��̣o�@�y}�u��>���k��(��~��jQ�"�����[�'�=�諣�hA|���o���q�ު�ޯ���`t�,�����g�%�Ũ�����+�"K�Zt�j��q�µ��&~?t�y�>T�i%����4�5�89$XZ1	(�ߥ�XWK�F>��ͽ�g���}��!��7��2�N�r�����Z�B��M�ֳ��5g���;
��¬t���,���O�2(��^ګ��;��v��}'2Tl�>~�Oћ�2�c��֯_��UZ���E*vO����^i���>�,z�ɇ(I��l�)�)����gl����)d� �!���	)�-��z��6n�T���"�wG�Ø����ӂ��)�aJ>�}��B�Fq��k>}2򜘾���كN1<G�5k�ݥ��Wو?�m#3;����@�<X�����.t�R�ˑ#z�{�ı��ޔ��,��8���1�$ͼ7WǻzǩW�����g%;>1?ϻ������� �'���@�]�o(��ψHS))O%�φbR&�ǳ�f�7G��Jvd:�O��'��P�Ի��$�'N؟;v��*��(��?V�u�d���W�Ż�_];5c��#4����<<V����'�#�����$�'�U���a�?��} �Ä���p}Sv�.M��5,�t��Y��92�a�j-�,ҷ"��w�� �������)l�����C�!b��q`h�V���;��%�>l�cӸ��Ů,JDM���s�ʳ}MD�G�ې5y���I}h��9-���=76���|���;���@wŀ:/{��`g^Ɔ/푆�j�a���G��Q�t8^��|BW,X�8�(l��cL��=L���`������p^����0��EzV�����<���n����~�[��뮈��7�q��m�ԳF������X ��*.S�>�+3˓⃏��QI�F�!��Vs