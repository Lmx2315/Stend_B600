XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��q�=�L��IK���T(�^D��d��γ5���!��7��O��W�s���~�ϝ��7�X^�f�W���{ϳ���1�l%�9��Y��L��r�%�J��2a�Z�&$|^(8�!���o�$���-�a��NP��F�l�q�D��`o��p�~<��皚yVI#��[�6�λM����FB�ŕ��~\�l����J�L�O�����5���Y��э~����sWҽHP��6�+˚��Gx�K���t�V�����Z0�H�p��O[�"|�"/��=6���/���H��iГm�+x��5�=g�tZJ��9������Ë�� )*~����ބ5q��b�}!�os�G+#K��$���Bz�-�h����`�c�6Љ��gr�k�ub2����B^�˧ш����ǈ�%��)t)��S�/F�e�Q�JpwʌaaD��V���h�P��
"2U����=9m��\m��#(	�&qO.i2��'yֆ����8�y2��t�$u�3�CI���B,��IjlY��@N~��f�'���c�ofi^�]"���6뾡���\��T^��<�:���ΟAڑz�P;^��**�i��k����As�fN*#H��*C�Έ{N��@7���1ȱ����^���:�d�]�v����;���N��������:�c%rfr�>լ��8�������6�aA����Ӿ|\�Ҝ��(��e�1��0*z�}Ȝ.�����,
�N�k�9��5HtXlxVHYEB    41c2     c40bF~��0�R@���r��B ��o�fm�}�}[��w��,�1�S�HN��j8x�_���$�}����cT@v�uO�6jf;�} �R/hKږ�P�M�8f�U��,g��"�
�
N�f2"����У�p������0�ŮSs(��q�V~�X�����K��*6)�4�"�?�&K���|�M�����[���b��a۞����[Ja�&N�ͪH�-U��v��h�x0<.p��P+m��N��%~��t�T7X�XM�aШ������'�jĊP���I��YG'�+�QU������J�]-hi�^�soT`���}m��TG���13E������YQ�� �rW����U�KN°l@���#ZB~J\K&�����A>�8$�G������s�#�(�a<�),��XL+3�&w.��,yn�35��b�nqj��6tr�j@{������v��߈5��ذ-P���s;O�b�(.v�imFO�b�Äj�I�~�m��~�|��I��5�	�x�߷S���7��I�'�J������E���T�����*��,~�<�Bh-�u��[�ϖ�-�����\���[���I<���>�P��q�.er"eG��|���h��b�KȊ�ݮz�8F��p��(��ɩkw@�\�-�9<qۨ���5��ʼǕW�<�9!i�4�"��xoJ����RvL{r�x"u��-;F�.f��,U�j�S�o�'�tu>�lkUi�D����yF&D2�)��\�l(��)�I5Hy��@y�Q?�cg�5���f��]��6*8fE�(�ES���W�>��;�Hx�FZ��7.Y$92A��E�6KN��.|M���|��[�[��P���@�:�\v�"���~?c5g�]�86F���8����#�՗an=�8�j��%,1�b�HSdߝ���.h�������ԓUt�_s�u �;$��HU���F0��4A�1E»��y����7����G��A�yZ�%���>��/E�"W�96r�5Ï1�U�@g�˘����}��hM�Ӓ��H�K��r�l)����ڦ�Xo��j�j�'D��FD�3�Z��{qh+�LOe�?vF���`4��USl�
P�LHp�_�7)j��2���M���H���\��I�LÌR�K��k�at{/Z����������#��d� ����E ���AY9w=�a�G]]�-�|y�Mg_�*rȏ�<ݶ!��O�b[NB^��kDE�=`��ϒ��:b��\��ab}��| �N��v۸��F�(�E;XC��R�:��i�*��j#�����[Fi��Zi����Q{/��漎d��A�>e�l�@Ⱥ+�2�ߪ��èfg��ܬ��$7[�Mx���ꍢ��^yoTǆ��"�������<�p�h��Օtēw�f����`�h���AH��='��^�Ϻ�x��y��Z�uW��h�I�@V��5�
���oË)���]=3tdi~ƞ`�]~�߯�⫡dv��r��ڼ:��X]#a�"y\ v�׌MS�S;ttk!ٞf��#yq�lV�/b�As�N��Le�\B����v9%~$��(��s0�ұ;+�J���=��B�#��n~�#!	9�fT�;�y�� 
���C��`I�D����Ƣ��yrĐ'�q��<���̓�\�w��P�	��$2�.���h=;������(�:�{�5�P܎�o	Jӝ�Ub�>}·���h���͸��r��tڔ��k�w|�2����.��fC �H]&�"�N0Q�Z�����+�F��xL���[�����K]*�O���_�9b_�X��ї`��g1[��_�p����É�ϪY���c�B�$�Q���:�#��k�Y��%x5"����`Y��+�Uv�sE��ilKsm�8Z��"��hxh#� s��&�m�A �O���_l�ي�:�\1V����p6� f�3���1�,�JD-���a�<��}r��yX(�Lt�BK)��t��~�E��:���ܔ?��\�`X��s,��2�:���Hv��G!i�v7�US�� ���B^��_z�91;��à�c1��`���3�آ��E>�I��o~�ɥX�,1Dn)wT1&�U&��c�]W�I�6ng��C�Q
`�'rrg���1 \Ro�ӗ>�\�� �>CF�/	�P�/�e�#�4ks��r[���O0GR���\K���ƃ��Ű�L��D�v=���M�`6��P�1��K��&u��-�:��UH���n�h�4��trL�E!�����I��4�[:�#]��iҥ�q�ɨw���.�͌���O~y�z`*>����y����f�UՂ�'����Y�ڻ�d�fl���4}�.nי֎�p�v1L/z��+�9R nm��`od�f�h���l-)ei�:�6/���=�?�L|�>b`��la��EӾY�P�)�UWSIĜ����Ǜ���9w� �M9s��*�PеsS")֎����I��)=vق{=���2�<f�B5�-h�^�S(qEd����b�S�� �'
��z?�z���������cE�lٽ>lZ| �R� ^��v�[7�A���C���o��гp����7����%�6��b�q�]�^6�p�R�����f�>#VV64O�ru�s��!�D#��_*�fM\��M���F��0n.��6���t�[�tN80�VP�C�H� 5�л(O�=��	�72�P�ٯEm)sќ��)�n�`].?�,�]�J��&��M�X�+�w�|����e�Ee��<��x�+�_h���9%s_a�_��օ
��������c,B�@�غz`����|�9�h�P����l�׉Sa~���З������8U�!!��a��~�� ��bk�5��o��{��C��Bց�u�:�[��>�P�U�+��%�kD�-�}`v��w:�w�v��!|[x�('���x/":��N��f�&�yi��7 f����B�h�X?�@�1s�2��1�o��N\�'c;Q�&v7�-d| L~�?�ߊ�^n��햊S��PR<Ae�ܔ