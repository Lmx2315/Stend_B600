XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��k��â�ćt���ч��
�v�,۫ӽ4�p�5���3�ȳ�jP+�w#�m��8�-_��� S|�*��>Y�X!�hL|���Ⱦc�f��c�_?Û��To�zOR����[,$˨^����0�5�G��6@q��^% �#�,c�5�	�L.о�� CRF��)T�Ǜ��ˮ$ж�وP6<+�y�2��6�*M����)3<.�I)Fek6�B�̭��KS�4��M�t`�3����^=<�yE��=�G���]Q�zV�N�avR�Xk��\�ZV-�Xu*����q�
���q��{�o&�� �3�;����>�iOߎWv�A�5�lV�	U����qD� ߭g��G�s>�	�!�m��b�`x�m6T^i�J`(}M�/�{l���T�J���L�Sp��f�[ĕ�z ���:����G���v�D�7��v�-���u�Cд>f�f��V�
�>B<����Ǫ��\+�~��j�^/��8³YFk�p�S��K�	�� ���I��jI�]1�e# �������5����[_8
�`�9>���$�D<I��(��*��������M��hHB�2y��ൺ({<O	��/o�m�a�����ixg9p�O����i������x�㊰�-;��3C4��H;&BΕ؍e��T�%.дE��"�ﻭՕq
��H�~���R��#�����Ѐ*��<���t�U@����x��=��ɫ�Ly�/P����c��XlxVHYEB    3e51     a10���}ԾtԵ�^��ʞ�x��MY��-�&Zl�|l���$"V�v�ބ��m��(Ʉ��p蘆�(��Z�B��l�0^�C�T\��ћ_�`tgf��3���I:s�Ǐ<�Q���^��{��
���J�#=�⇾�(����m�e�E&c�`�mF�M���d�!�:4by���P�u��[��I�e�j )�G��!�uC�ˎ^b��6���;�6�j"�9���3����ܽ;?/��	ٹu��}(������j�M������بQ/�ȭur��>����;[��V�h����O��l�aKm�<NC$8Za���x6�����)�`�O�//��6�4Fי�*�Q�ݲJXv�r}��8�q�	%FW�	8i?/�6.EP�� �����������I�Q�GH~��V���ѭF��C@ҽ���F��\=��^"��MxrC��c�z�x�"�1Q�&4eA��?�#�O�����ͧ�a|��5v[>�����u �fPy��+Z��fi�jE���6E��I�~���΂�=���]�l�B/B���t$ݰ����Pi�j�4WdW�gk�|���U�f\h<����/4bD
���I(v�k�I��#��PR�Eo�*��a��y�Ù��[Wt����q1��5.���u��N��$1���P,�D4ů�{�'��J������l�����A�쪭4i+��]���ۆ,�nT6�]�+�k9�e��F�	��r"��������D>����8�n�n]��S�,(�m��N�3���A
�^�b����M֛��2�5��V3#	[8�$���W�0���6\�cX�V�G�]8�S�%V���)��V�t���#�s�8�k�8���Z]ﾴ��F��Z�����*�:�W��ą�?	*_c�塤�=)cL�DR���d����X	��	sq� �%��"��j�6���yg�N��Ց������ɅR[���� 	�L���Q'�;��z���5�D�{���n���0D�{0�AOe	�rWc��6~�1rfJHN���5�l\˚pU�n)1����Y��$�|�g�jee�^�["�c��,�*[�,��X�d��6Z�7j0|qo�i) �k1���oO.����#��8	?�SX�=dU�,uΆ?̡����O(|f��d�*� i�MI!�d4�lʖj�l��"!����}�"�R]�b�3��xR�O��������@w�ޫ_U8u���	&Z��G!���ӑ��%��4��_?�7yӫ����\Z�t�0x�1i����t���?BtI��c��>������uj\��v"G0kN������r�ð�0^�hL�aW���?N⾷`��-��'�沩,I�kܯ��uEi���b�4B��(�}�?�:BX�ٜ� upc�Q�.0�z���T��d�
}�ER�/p�k�2˚�5!D�A�>�m�@�EB���{�F��P�,k4R*��:y��!������l�yʾ�+q�T�2{i���Y��L��uH�Z��,�08ݻ(ç%�,
6�=��>�H۬(*��cv
LW���ZQӦip�n|v�	[�4�#"�בL�.ʤ@W��5"��qd�m�0!�1E:ݱ׫�	�������1'�� t��ᰰ���q=_|9M#��=@��XJXRҬ:Rt�웪=�BG������з*�%4lqX�?�Ϗe�7����w�+ل/�ؓ�(N�`�M�~:"4vH�&
)�u�0��4�����mP�!C?�� #�1,�D����RX_�<���:]g�$�Y8��*D�E
Q����^12y�Ə��>�����q�l�'[ttڄ?Rѐ��� Wq%�#H|�&$�����xT�b�$=�c�S�����(�F��v\v�L�}�v̋����ହ}y�scK���TO���ii�U5*��p�(��F�])[�O��x\9#�8�ش����z��3��&�׆d0U|P�\�Gb�0Q��1�-��LJ+���eOU���ӡl�~���9 �Z��Zl������Y�4&�2$W�t��X��&��!��%n��ªێq�	��C�m�၁�ex�T4�*5%ό�-���#�g^vk�\����?�3|㛟��j�!O�OL���垬:}H&��0�#ذ�@�~�Q�=���gP�ۦ<�)�-]���\��9�5�6�-8�
����ݱ�Mn��J��	d�VIT��@r���X	񭍴/o#�f7����U1���Mr|ٯ/���VB��0Q����
]�3�n�Vn"l.���3L|;�`�?��G<.���?Ȗ��S���Wzԃ�$g�iԯ[�u�)�����:��L.�n\��L,��z�>Fr�zPv''CuP,�^@����(�]�MF}�-�����BgO+��Q&#���}	 �!H۾�:��Z�!�ޮM1/ˮOj3���S��x��ӣ��zB�̭is����� A*���g)QeEg
\\���X�}Fق@	�^5��L/��>�ԡ�*W=}\I1��b�p�*0�	RH��Y`�Ls�h���d�p