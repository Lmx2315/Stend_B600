XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��]��b�\�Yeb&A��_#������'n�C�gu)6���J1LJ�	�0J�A~�s�R��l��{(���,x���lj�E�����t/yd��=;`?{g��EU�幫?I��˦MX�:�����:S���M((Z�$X�|D$��e��_����48'1/Ӂ�j��+�=�j�P�t�-��*~�>l"���A��#��W@����sƗ~�Z���$ζ�	�� �ٺ7i0\5��8�ބ��w�uͽ����P.�jE���u$l#k�y3�Z�s��ԚtZ�wQ����.�"5S]���ԧۑ��e����4겣	X���]D�E�+��^F.��̕12�0:�|�a��Qja�SF��̥��ȥ��+�:����/{�@d��M=R��m��[�K$��h��ɝ�9����V��%���3�"z��%.>�6�L>�q�B�S��:I����0�p
��,Ţ}��j�\�92�4��x���2 8t�.n�����P�!;���?��'1H�F�J/��B��s&�N��|�P$J��%EG�8\���k$[Q���[+�4,�9fF�?&�yF��Aͽq_��	b�^�,�&S�j�Ƕ�p��}�θ��I�SK�ȭ�G��/�hIP�=<�h�W�!x��%�fv�,=;؝�e������S"9;�$k���i�C�MZ2�	�"���8XN\Cw�H0j!��;��%���4����f�S����:�l�X��V��%^��C��u,+��uXlxVHYEB    2902     a40ҳ�Q@��_o�ucXOR��v6Pu��&�����(�����s���JP��?�3�\
[(�E��,&Z�^�=�w=��n 2ib������i\vt��.��|,,�|��/lXV�2��ܘ�8\�R�1=�u��Ku�E�;�8Q���b[�P�3I�ҽȇ��H�Yu5(�`ۙ(�8�5v���_c�-��sPl(fC��8^��:�E#6��t2��Y�ʷ�����nLOPJ?@�	��ù˵�m!v��H�9���-m�Ά�Ts�̀�DbۍT�{�n=��8���=�Cp�Ѽ�Z����נҬWߝ���c	_cl�E7N)�8_LB����������±���<� t+k��ڏh��3�S�P���+ܔI��V�)��9��+��Uy�#�(K�p.I
����j0[�s_�b���'j[�2qD��2�V̅h��������d]D���#�/9H�$]u��ȑ+P�y
N���&K��bc�+D�}�7B!_�]�V{N=p��Gx�\TA�nTJ�PA	�9r3��OL��:����ެ��%�(XhB�o���tѼF�ƒ�Ig2�$��y\�Z�83��Dp(ͥO^Y�M�:���P1����#�4{�����y���?��P����'�6�8��l�E`��P���0��w%����;w���?�l��t�]��#�����|3x�5�`�dTb�6�(kϴ���I�@�b�[&T�p>\#C*��ֵD���߼c�RmսO�I�U�= �%o�ZGA�ZWm��1B_4�����������ˌ[�:N�1��&Y��]�X�Gii*�%.����_[v�{�~jNٯ�&:\$�yEڕY���N��/(6�6"=���%��!#F�uM2�����>C�j���}��|��{��e'����Ea�^�Ƹb1�����:��WF�XHn6F\+�w�g#s��c��hgK�T`��Q���r5?8	��ۓ4_*�V��)v9��q�I-�d�n6^�A�����o18���=��\�Rq�T{�O/���a�\�	rğ��T�@�ޝq��s�#*y��������%}���С�yk�f����t0�����t.��А��H��~[nS5 �?����}a�1.�V�~��c5qLHL�31��P�Y�N����)����?Kk�0o��7n\�d����4����4"!���a��;D���t�~����.A�N�V���d����(l�F�w�3ێ��>Fia�U8�zY��$+�c�'+a5#j�)�!!$�\��bY�K��3K��g#��+0`��%d�4���c�k��?�+<��>���.�b�eX��s��ɬ��]�V`:O�?���a�}5?B��)a
������*=M}�^�zi��%n��S��e������ZJ�:+���D�;�<B�-�A�{|�?B�0˝�8:�z
�Z��P?J��ظ�7+fAǤ��"�< ��G�K�x�|Bw�D��q�2�6!�EXV ��!��@�R/�_z�]��w<"s�t����ь�p�`WK6pzh�	�sD����<.�,Z&>�)�$�ϸ��6Fʠ"2=�M���@G��³��z���+VU��!#
��A|�z�_�q`�lLa�-�[����	mj]�������T7ē6���31������ɻۣ��vͪ��;ױ^`f�׈9)j�w뵏��OjζI����ܫ'��7�sX��x�t��8�
==G�Z)��ÚX�ŅRaAw`x���T	�J��P&b���G/l�W��5����땋Sl2n�#��e�{�P�;o�������vU���v�f����1�]^5�p�y|&'�
�<����<�Yf��cy_+_8����(	�
pI����G�1\�\��nM�Q��u7`���e�(��+�ڶ�����V�3#_q���9�ߊ��F2 �e[��o�/a�~�'g*�7.ch���DTc��7\�͒�s�q� ��X����'����4Cb��2����.�~���}PQޞ���Z�����wf�cI��վ�4
gp�)�HƩd�B�^̇���wh�����=z��?C֒�������C�I�\����(�!$L%Isܛ�u��x����{���Қ`��a4]��r	��.Vqb��o�l�-�ٔi-t�����=T������˝�~\"��Qܷ��P$�T�w&��y��{�y�㮷9�V�m�!E�9�J��*�&�찿p� 3Pc����,���X�m ��*��_S�\�h&�(m �n������l�m�c!�������7�ش=A1��q(��[��!���_`^�N0%�XF��A-cW���Ao^��r�)��tv���u��m�� ����Ka�Os���༘�t��/�K��k�3��G_ii��T;W��y�J�韲_�0myT����ZSs���H��/p~Z�~�����}�e��~{��'y��<�8h��I��Q#��������n��"Y�0�q�9F�VÖ�Vr��R�^=F�]w��R��K#y�Σ��Hӊ�)Q},��_x"$�Oa	�9G�}yB�