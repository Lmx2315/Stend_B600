XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����ZN.�W�|�PQ{EZ�F44I�'`�����2���|r���������OQ�&���XǪh���Ƽ�M��^,���iG"*��O��fE{�Qt��R�?uB��=�\�EOL6�l����0|�����O�L7�dJ����v���������gTR�{8J6�n�s��y�df��`I�r��6������o�r+G� �����=�I�+hC���QQ��*�7�TZnKk������	��H������M��\d��1��t�3�������?��E}�|��2o�ōu��0���(:P����K�yv��=�C��urD*���U�*}j�T*����A>ߒ�\�fW�i8 md-T^Ρy��D�R�q�`�z�#l׮���s4����Hϯ���G8-��<%��H��m�i��t�ऽ�C�Fs6-P=�r4F�r�i��<�&9i3�����,(j�z�Cɣ��s\xӝ��j���^W��L�����3){i _=K�ty���3};tߗ�̜��~Q��p�!.�h�#GL�غ �i < �z�'4������{GU�� �ٱ!�bJ�N~ߨ�CA���o�2&NV������iF���l�;d�x���+����sN��`�vrA�@�@#�gt@ѐ��Z{����|Z��D���:�7'!�	Z��W�`��9��|_�Gb
:���_B�����4�� @�XLP͎J2��ea�� !|��4�F��zU�T<
WE��x�p(��XlxVHYEB    2864     8d0-���Q/����ќpG
��u�ɒ``ⴡγ�fB���e�8�e{#����\�����F�$d�e�wzL 3{���Ѷ�Ʌ?%�rї��|�B@����_�jp"���қ�ɜ���N�g���08��qB#;8I�4�6=�y�I7�?U��,&Fn&��*C��y�v(M�_��jET��T�k��ެ�k0��_�%�>�����-�QH3�����K��=��nP8���r���Vyjntܐ�Ef�nk�r,D��j�G(1M&Z,��k���yw=�DHD�V���K����6�5qiKa�{����a1�#��A� �i�K�l#�@�j�����8�+��/!����`�C٦��ls ��M���Y׃)�p:{ig��ub�&���$�E�@^Fxr���LaYi�p2_x
ęMS4��DW�TK�n���c��D��w��&ֽ�q{L�`eʅ�{+�J�\�H�0�����6
�G�u�C�!����Ckߊ��W7�</R��闕�$B!|Jq��o�����6��W)��d�0gU�p/b����$���ro���Q�وdFXD7�� A�#����۞+����U���X�뚥�ݿ ���V˱������Ԛ��;x2�BK�V@N���1���Ԁ�a�d�'����V�Cor��g�,Q�(� �!�9_(haH4Ĵ�rjRJ�c�#Y��<��}<�����&Y�Z^ȚL���Re��T����[{����{I�P�]B�-N�߼����6��<��!W�c��6�v�U�T�����/�@���GG�t5 z1"^�o�G����?D�P�M�C�Z���TΤ
F�P���;T"��E�k�؞Ě��L�R�K����ߑ�U�g=�8�$��s��UU��elw�*t�z��ޜ���e	�>�wOU��.YV��r��7���8��YB�%G����v�3��ڜ�1�����B�kQ�V�$���=��?}_��2�j�>��@�v��������P "S�bP�2�� ��:�~ɝIF��4�%��5X�n�xSYA�2���!r�:��pU�.�0�Qx�1�����h\FWrJ��b��y�U"�1��5�X�X�s�k�vL���x�?�:�૸��Ծ�Q6$����b�ǞbF��V���}�� <:�fe�{��%�mc�Sɨ��!FV��o��S��%7�e�{]ʻV�&��$�`�F������G!܊�[]]�릅�{��Ay�\?`iW����G5}�&��P���4�WiJMZ w2|�U�GXu��c����YQs&Ǟ˻r
�Q��h�x���p��N �c����X���1��H[��(�M~����9Z��be1��˗����+�؇_Vr��A�,�}�e69Iy�q~�I']7���n��Ϊu˕:������-�HZQ>^Ԣ��E[Ϋ������F�ъ���%�x<��Zs�|1KF�θ�S��@�1^���7�6�����R	:s��V�z���JS��w�QH���:v&��	t�(�$P�"�S�4��s�3��t������D=]��y�������n�8�*�$�E$b9,uo��l�%��92R"CrdĿD��vWb%a�[��k�xs�=N�nt�h*�n�D�07&�|I�<�|�t�d�@�j�|��x�W�)GpG���i�J��(��
���P^z��n�,+���l�Ԕሗi�3�i�nR�gB��M<s�\5���<�[xz���U'�M@	���n}�����l|װ��N�FR�آ��0
$�j�R�}*���=Q���N`X���k�xN���.� %|V��m5
���Ia?C�$0G<�˛^��_��\�c�v��n�,XO�&�߽��)�̲��%�e���hL��=T��$�WK���*79A-Ȏ�fa���A��{��b�B��n�8�D�mߝ��l��0�*��VR��Dn	,�P�B����xA�Pg8K �{��v ��L��4�`$�M-2ɨm��_z��.�A�5�{St���5��Z�A�uO5�O�F�7��T[�/�Z�*���sa����š[�駘^Mդ9zE"��;:�';H�f$��	Pu�'��X��K.�Z��i^�>��b��isJNV�T����رU '�3�,�8현i���Aŋ��c��뒪�g|y2s���y ��b`��N~