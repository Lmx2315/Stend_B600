XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����y���R}��]Fk��݃��y�����s��Pa���W�\�����6
eC���_��3MJ\�щ��9W;ι��cG��<�C� "��e�'�����49���4	!kй=��#�F�9H)q�c/mM��fۘ�gC��yk�7D����C�I��W⍥d.
�>g�1д�S�����s��nFi@���1��]�V`��=�<���-�6�\p���\,�8'�Z6,��6���H�Y����!	ї�B��#"ʇ�q2uLQ���o�ie$����F�ϓP��c�̂I����K�d��}��T��)�����)�3Ȏi���gb��F7u7Ep���E�w�3f�L}7{<�z��(ΦO�u�{(蠓���e<s��-p�������|��S���u;V�v���(3Tm��aM���X&��4+$�y� k�0��9�MBGUMq�b�͢�	xFʹ���;��8����E��N�v�}i�p�|����t��*��N�ˁ�M0u��&a[��q{"��VX����k���g�fX��s��ل��|���5!����FoW���s������,�8;���-���Y#J7�J�����]Dg��������rW�'[
��Ղ��4ea]���!�;o��W���H�Π�"���q>����7� )U���}(��S���N3�t?��V��%�5��������Ex��@n���MT�$�A@��3��=2Ez��@b��)5.�5q�^�[���h݇5���4E�T�謟d�xaXlxVHYEB     b05     370T^�C>�[ih��݄�W�9\WboٽgӐ�~�Y�f�KJ��`�yn�&C؟�ÛZ�5�N�J��Fn���L����ΫߛnP�o�I�}3)
Ϋ�S�
A�[�J�]%�V�`��e#|�p��*�Z9o��RbOC��%�'��А�oX��C.�"b�8L��+��(hWYu]����S<��\L�)�F:�n�}[^v/�wSԦ�ڔ�s��X�I��5Dw�m��d`GU(6k��(9#����yń2rWKOU�ֳ�T���&���$��Q�}��}��G�x��^@IB!GC�7����W+�0	ڙ���ϧ�ÿ�����NG�v	L��W?d�k��)s���R$-/��SĺR*���k��î�Ed���p;a�!���V]�������c��ـ:3�;���O�Q�{���pxH�Uѕ�$O��לX��ҞG_�_@�F~^l��DWƐn�%uj��v �����EK�Q�X|@:+B*ǂJ�n�Z�(�	������e�q$�-̕����;f>H��v���'i���Z���&��9s����Em�cTڹ�EK�	��FS/_�u��]�R�>EU��1��-B������?�?��cm7lDX�-C73��Zt���P��ns��G�<b��	!��hS�')C6�K���SZV�9�}�$'��C[E�&�v�� Q�Ϗ�Eڝx5>�6GMNr�K�kjnUI���$A't�\$�[�_�!� э�1�AO���F[�ե�O�QQ��=o
���(tB��n&15<�'b#[F��
��澍����+���<���J�n��p<�Tro;��`˚s��k, ��)x=�f[�:u��V&1h|a� �J���7�cW����