XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��E�]��1d5�iy�KP<��!��;\�'i�����99���۵̔J.#����jۈ���
��r@#��q9��m���0��;!�w�=㧻�j��\T�>u�������4��X���W�+�T�~Y���5�+�x
E��K�m﹢��D�/F�(�44��X~ ���I�T#���%j��x�B�^��ʴ"����]�$�EW�A!�!�%'�0ã�J+�~ޘ\RC��N�_ì;N����$~z�α��f�؎':������)����X�-}��װX�ʫ��nx1)��R�'f��@�I���u\�q;���7�E���a�=��'y�e��H��=���l8�5�����V�R�g3Z�;m/��G�ɝaLb;�o�M�G�D�(�B�~�?����f\�@�l%�R�����&Ъ� eN��K�=� �+N��0��tز�B��P2I�0|K�RҗbS�qrs���P� �B��i��N��G���V�fn���w���Q^�1�WU&���>|���H%��.(�1���s8cf!O��bE���1c��U�����
ݽ�K�U9ޅ��3���[�E�1�@��p���8p�fǔ���=�2�dK�jmk&��� T�k�Mc�����J0s�����pH#���r�\�\��=���-m��fm�|��@�,V�X����j����R��:� ��/�eaa�[�ߤ���[��13ʙ
����!w~��!�}��ЃG��n .R�E}XlxVHYEB     730     2e0P��%1�}�W�d��k�x�b����4*{���G*�������-�B�s��z�i^������E�_Cp��O���}��x�J�]+����н�u�v(C��9�yb����L8Ӿ�T���`��3
�~3vR
^�h�(7��/��h&qli"��Ǒ�Z����P;#��-=�[�i��@%�֦JO�a�jhbPdh�q'I 1�����6����5����j��X������a�4�@z���e+o������Bd��Bߡ��M�wH#�=�h̟ �����=��o��7��l*��I����">9�yť���������t�����k㨒�ȩ������jp���F��W�i�\�g
=�:t��D�aK_�����&^��	����ڽ/\Tٴ�b�Zڣ����@A���%k�6�g+��e�,�f�{S/NHO����zW�aq����<�����e��M�i �Vy��G'�uR�&#�������W�ϫ6���.�J�<�;\#�>;�FKV��Z�qf�^=�A��v�)�ך�Oiߒ���q�-K$�Hs���U�:��0A�t0�m���Ʈ.n���u������e��������Gf݉5����2��1�om��/Z��X�Rq>isS>�h=߽E�����=���N���Z�$�y,p�񕥈s5�>u?��mJ�؉� 顏,���h^���xKj�n�A