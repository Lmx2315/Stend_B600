XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���-��l�\��m]��<�vr+ 6�C���9�x�����fw� ��X� üx����g�gueJO&��W�O���:�eA�׼�=�"�v���;��&/��y��C�:=�5W�$��a�yMMӟf�XWme.��՘7K=��z�x�����1��ݕ��`��i����gU�/2���E�>D">���ሳ�y6@7G!X�<dЦ���4��F���o�(5�)�DC�$�=��&�u�'  �V�!��Y�bBc���̾��xs���jB���m��I��C)_Ta��w�T3A��+����<D��
�5�͈A�����������ͶXY�F�sg�f�CɩC��h��'zZ�BW��Q�,»�_�cӼA����x������3�UX�5�����X!�Y���x��Û_������>S�z�:�^Q`�]HyQ�O5�~�6�''��*�	���1u=I���{�Z9�Őzn�>�h�B��3��[�X(�	_:���585���:�0%�62���t���XA>1̍j�a �;֊�Րt�ث��E���Y�2���A@�`�*E$ؚ��P%�Z��V\HE�9��zJDj�=k��L=q{<��0 q��ouO��y�-��(��ϯ�uHO/���ǖ�`|��]���G�t�6���A"��˸Ԛ6/<���$�J�\��>eI��m5��|'x%`���[2��+�u�����e4�o��b�l��w�x[�4>ٝⴏ�8��oλ4�=1��XlxVHYEB    152e     580Ć��kݩ�,��O\݈fWd�N��j?���XJ=q�ժz�x��}�pj�YԟӢ�/.���n�)]�j�����c3�����]�ao�A�Q��Y� �@�m���e���R8m���l��N��:�81����X�B��j�ElJ���ƹh�R`��Ⱦ��A�k`|����H�``c�P�����Qq�08��2C	a�
���E���heu�pOo�L�4v~㋮�6�\��%X�mbj��v��rA������P~
E�pM�h��Յ?���[�EiQ$r��������J����F��N�ZHi�o�aI(��G"��'��T�YU��@z��#�i��a^qXz���;��h_���͹�ƕvOI��dm�����X\�C������E7�v��Rq�7l�ר1����s�6q�H,����U��(QTy��h�>f2k����Fe;\73�sg��c!x�2�/�p��.f�{a�/�)�9�fr������F$�/���PR4�pZ��l�u��Yu��1�J +ՐƎ'jy)#ű�^�f	:s������~���ya����OH�t��L��A:+��~��[��m�س;�	ϊn�}_�����k����#}(�.���әi������mG�w6P��p�;@��kqۅi�輪ȗl�?�M<��/ g]:%�۬�Ԅ�Dݺ��Uӷ�0��ߝ3�b�@��dУM��>5]��A�7vP�)
A2\�$�����С��H9���~�x=�M��S�����mn?n�p�Y-�^��8cd���,8Z3���|�X B	Y4̴�9��&"o0�� 1��Oᖾ[��m��Z���f"��P�0"	���o�4���w֑��P��%�/�
�7m�6�GI'kA�1ܠ�F|�e"~H)جl�Kg�"�0�uR�gb��*�P��6 Q��B�S�OX�Êp���~c��~1���-��F�~�����T}��i�p�?*0���P��Z>v��x��U~T�S���ɊTz�E�	�o�.Z�޻��{%]r{{���g�-�)]��m^�l�.β���z"�?1��8&lU9G��Y{��5�`y��=Ch�Y���p����i�T�����r�[�F=Ռ�u=>�+u�z� j�.�+���|g��T�#%y�X@#�w��+��W"3%UI�ЋD�L=�� ��<7�a�Eq�/v��E�C���9[+�xk�Z�!b�o���zh3P�~H��(}L��I^Ä���gS��D��C��X��ۼV���߈�)���čû�ࠂ�n4��*��r���//v��SxyG8m�VZN�BV�q�X�Pӗ��� ok 3��P�����NGW]�:��������=cG��Z