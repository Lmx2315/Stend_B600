XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����f����9<��j@���)J�����
M_@�-o�W�՛xSe�ݠ�(� ��JԾ�HYh���3Y���5O�W(�}G�&��DCC`���3fk�]�٦�`�J��A��(FW~�A��iгS��  )��n���A$�ţ:���>.�SH���͝����6�(�k�Pۢ�!�xt���
`�E2��C.��&>7zW��0E�G�Q]���1��w�)��G����^�fLb�N�@T��,x���1��Zg+pܘ��=�mj�yIK�"���7#[!
u�Ã�e�5d�m���uGd|��#"��!�	���'�U�O��� ;:Em0���@��F��ih�ӕL�4���|8Lg3���!�����jjk^��J�G�0ޱ�x�2X\����6���\�^>��0;�ꫤ�������W��yN'�h��!�ݪ�"��#��(��,[��gj�W���U+Sa<M�2��5ʭ*��]O2�͊�&�E`d�B���cb[��I���&�$�Į����#i����båe.���6_3\g}�5<�(2�rJ�����'����f�����;ꓒNF����J^�㉲�t�6��R���e�l�t��z��g���7�U�jٴ�wRkk�趻��������Ai�C�Od�j�)^��weD3.:�/%�>$�kW9y<>W01R9';��y[X8É�V��ܲbE�>�� �/{�擑��~Eq���_�ȉ�?��}6�/$&��{���qďl݌2.۽XlxVHYEB    27ed     8d0:�ߺ�#��|*�iV�y��z�U�j�$�}��٤y󁝻Y�w/��v���u��n�׿�jɊ?���D�-ꊟ�	���Yӈ�vv6��]�L����Y�hz#4��Buq��}�}<���@�m|��v��y�˅6ɷ����6$�/��<��4^u{!d�֖��#Ϻ��d���H��I<^7I��m]{����现+"�ifHϪ������-$�ig�f�LJnk܉<4�۸?z�ZgHo�hu)�	 P4��pQIm�ܖA��޴W9�g��/.�\eK��[���<*`�A�*h��W�y+���+>����$�?��V�i����}�ڤ1��Bf:�̈�H4��m]B�+5���
s �ۙ��{BV&VK$���Rh��;S�q�#�w&�aי�U�����A)�tb���}D%���	�������(�qf�Y#�t8\H7�:힠AL��B�<��a
�(�UB ��ߘ_��n�^���0�}c���l!����3è2p���eq�
��&����B�4i)M�N��R�A�[AȦHP�l��-PR�~�/�<=�{�#�1~�GGp¹fi5Bw��y�� s�B��/�{d�g�,�7�W�ß�Y�3��#	ڕ�����8`���;2��&ꨰ�1ٻ
�v2�È��O�8�	�� �	y-Sd|�1z����6���0�i��<	L��ڜD���Ҭ7�4u��#�����R&���An����L��6�p*V�9R�3OF:���gr���/*����-�l���_l�Q﫱p�'�]q6].��ڭ��=b���py�P�x � �@��%��d�E
Br�>�G��$��#�*#��J���N��Dë����Us�fF��0q:aGd�xv6īܸ?w���h #Cnx���_�1e��*�	BV��H��e
�7���UzP�9����mi[�or�U�O�_q���$.z��BQ��5�sY��Ocs�G&�d����?�����u"�x{�O_������2f���BG�>� :rf� m,����أ5`���<��W	�Ű���x5�v��Ā�����s����sg�4�Vt+��M�ʩ�d<&NB�\���T���(O��a`�!����G�9Z=�[Mj��.lK
n_��
3���W��������?�U������g���
�v딒Z��V�ז(/$��[Ue�ּ�.e���^B�a�Y ��I�=ѝ��w�>�.�\�1^;}J��V��!w�G2�k]��޵�	����=��"6��N������s��9}�� ����XJ�TF�UY�=_�������t~����!'*a�ʞuU̕���'�?Û {��ѥ��?�X;V#�|������Ue�X��\�74�2|I����f.�f��?�7��z�A�Yf<��礽`?�At�(��Ht��{��[��w��'2	F�ES�&g���QP�Ei���h��ą���5V&�Z.j��ד .�S]���*��
����S�u,١}��E���5���t}�T��"� ӿ�[�f�Q8���ŋS=O����3�V�ְp\�6�������Ԫ�.��;:H�[���%OOj[�]gä^�3�+A���=x#��Z����f�m��xJ%��J�|�.��;0�4�J��Ä� \O����2Xߍ�N���O� ��p�e�7d���Y�~;%?G�1	��s��U�n�܏�&�?݄����ĦC��R���)EZN�/���Ya靖��8r�m�
��1�X���&�a��n.ce��_`���:?Pp6��3�f��q�&a�g�!7�X^��#!������N
��N�$�pĎ	��[<�er�m��,B�ix�߮�IFVP�n��Bs�I]?ȐI�-@��X�1qۤ�e���e��d����Ѽ�f��/�]<�1��E9D�e�4UH�l#��?�C�ϸ�(�8�ɾ^��P���;I��z985	���3�!��|.�(AS�~.��x�6{��Nz��uT��|V~O���|�Y�@��D���ë*@9�l����re��{�b����//���A���v���,�3�щ�,�DI�g{Շm��6I��x��A���C��9QԸ7]eS)Ѩ[1�H��b��������^쐥K�j�M��a����!MYU�[B���[2.8����nu(�^�m�#2����"���y]{>�b�PL� ń}1��� b��=�l��9'�Z