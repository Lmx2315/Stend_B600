XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��X�e�6�m����%L;�_�:I�+��8�8gA-Q�K�]s���߀2��d�F'��H�~Y��l��`B�0َ�0����>zp`��K���0��Gݫ�BǤ4B�T�j\.��\K�b������9��>!Ѭ_�N���y͍9�p�stvm�Z��r�,Կx�&��.{��#QA~��9u�p����j��D�%ߤz�����_Q�y�4�EG6�@��I �KOp;O��UM#$ �H�,d1m]��/S@|	3*�^ʇ���Lx6�Zu$�����V5��r��m�h!�B'�t/j+�Mk�_DG9�#��*l�ѓ(��M�D:�%z�F,��ҳkF�����Kk-���/�C��R��F��:Z@�DJB�y�@����8?m�Z�m@qR.��M`~�J�dy�u��!�<4W��������;��,���g���A��7uwU?�D�M	A����TC�O�{߮����?t`���xi�:OV��9�E��$5h����q�N�xY@h���f��|��5�e��;�4\��<��zK�mҸ����bѬl�m���S���X�����Q�\�?��Z��MI��p�E�h�nWF +��K�ή�z�����N/��P!d���IpKi�_6�u��Y9ş�]�I�0{�XfO^�}���U�Fc`����PQpBm��l)�̀Al�����������W'����)�3��߹�f���[��D/�@{�q���&�<��*����`J���Q��z�\I�XlxVHYEB     a4b     370G�ED�|�I0#M0��@�ǘ�=��!?��桑�j�� �(8��`=#��9��A�A��kJE�ONb�\�ն�c(��aDs��G�u�MZ���3|���A�6��ܧ���);�[� �S5��zY)�J�T�nx,;Q^�&F|�:^w�r�b����A�=� ���l��%�;�譀*�QH�C8�0���g���.��ǖNlM��9v~�@�w�	i��;�T3ױO��ش����D��s�qU�w��x��看�`+��Z}eR�s�����1,猠ƴu=�D��uJ �͑V�|�,�xs�����/Sz���)���W-��i��lb��Ԥ;��ug���C	��2��OVw�r�1��mV�ɠe=������-�;���P�P���ɂ�c/ŎN�hOв?��9�DvI���cQs]�eg��yBk����(Sècؖ-�T��-�p�b�\X!Y��E��6<�eW����2�����6# ]Ъ�K��/�2����b�G����l �u�d6H��O�Mz��������h��
�����]*�c*�ç�'"���%zz3q�`"�d��L�a�{��t���C=S<��߳�<_Wg�uX�M_��E�!�:�q��F�P#����~4Ns��'F�SE@�Uk���0P�L}-&B�E��3���}����3[R��]�U	�d�k�81%9��h���d�ݝ9�����&���v�0Z���-���Sg��������;i	������@��ޭ��ź=����8?�w����l}\��n߈K�4q�����`���(m��q"���<�_i���CmЪ7�����&�[9��MH��^���v�'si�q��B7N��f