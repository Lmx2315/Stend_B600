XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��D�xw)N����
�_K�m�6`�)��1���7�
��cxx�5Z(q�=�7�q�:�w5b6F܇(m+�Es��v5������끹g�������3R����m
���+Ɔh�A�A_�#w��l�8�ɞ��?c.
_pmt�l�U8ņ�.���<��m���Ge.Э�W���]�P
���t����ai�`���缋 �iR�"n�f'86�.�G&�Z,1�Cx�z��/}d���q���!]jO�.>۳~_R�9%�_������v�6�LNd5)8H٬�{Yګ���ϻ�鳺؃/�gB�Q���tVP֦lW�@W0A�g�9�Hi�^��?#�=�'�a�`��i%4��Bx�٪��C�����bv��Ovb��:�{��6F��#q�y�f��z۹�}^ ���'��Jx�s��^�э��z��%�>��\9�7%_�Ȍ ;�ǎ��u��x��4�_�ET�,�BY�t_�>:�f��LN�4��a�iHkO6>E�i��
���?�m`�Z�x>��Г��G�'Z̮�Gky9N!��y5��!H/9@���q��4�Q��^�X$�����%�:H'�g��{�,�w&���� ����J/��F�+���(��$R�H��q�@���Qsʰ��O}m�Іɧw���=Q]@�d	Ѳ-ei�l���K�)t�L�%�l4��z��Yj�T�?*�,�dn����G3���z���0�"J^��v����73���6�b=��Z�mXlxVHYEB    cc3b    16b0�$�ΉFZ�<�I�\
]zp7*�s-�t�����q�o��ٽ�A;��a�r��WȷĹR��#��|1cċ�;C�8
8�I�'�_�f`�$sJQD\�%ŕT$Bp���Y��	f����U��MnO� ���h�����Ƶ�����q�Z�?��f����u���q�+r�Z�|�{Ͷ�����$�<�����#�ԑڜ���pb�(P�A�W�%��_]#êG'٨������O��rV]��4���;��,D�k�A��?������H���?%�&"�ǰ��{CUNl5g���Eɣ�¾��MC��5����ra�O9C\�	���ܜ�w2u|��N��eM��>�j�_{��3�Ԩ�>��G]L��.���'!N �-��?\2�>p,�|b>d�%��{W������M8Vekj]�,�v�f֘���f&�b���z貝���#���2w� �ˉ�p�VK$;�VzĤ�7b'𡦴��v>�Y�Odt1��|ES�+�fO����w"����3���t>;�:��Sw�;����:*��P16�^�HB�o�[.W����A�k���z�,�Y��׌���A��!���;]0mJ8	��}��3��4rl]��p��������Na2��Q����%p�|�g�`�q�A�k#a@�D�G��D	j�� �f'_�𯯬��@�na$�H���5��vy=t���\�����p�_Mi�>g��؅��A������1�_�V����u�$�AjGǾM�Y����4��g��W�AX`�H��A��udd���ʷ��M�*쇷�ѫ�\�Kz�e��uԽ��$�ʤڿ��<�;+ߓ�i�wr(�8D�C@��'(��^(a/J^�0�%���D�p����ib�<5B��g5����@�t޵#۩�tLT^�噘���+��]�{D@�f��&$��W��2�m�� xe	���jt��vEtB�'յe�����b�O��fn��+Y���\>��v&�P�ohfU�1u�-�nI"C%
 �+i:�L���0�-?�7|XJX��y������4�tŤm���џq����2SBwE�9�QWV�I}� ژ<���)��J��\�xH��-�Vz�����Q���[�;xp��1��[�.�A��!����NchPn&Q�KgX�8t+m�n3a�a�L@�M*���yR�$���!b�x��自��(]�A"|�� �o���L&F��~1��[��!����p/�;)��"8��a�KȬ�����	�85lX={��ǵ5LZD�٠�˨>�;��߹~s5ҧ�x�bvbO��'c�6b��O�����i����|ccT��x�������������x!�F�5��a��u��"YS��<ׁk}�5��ߧLe�N ��C�z���1��,���a�GM��^ ����P�$�᱋�4�SXS6/q��X�&���v�MB����3�c/��G��g�^�=�C	�-=o�5���28���]��%��J������1�بTm��sx*#� �Ɋ��f�)W�c>:��7L`|��ۇ�P#�7���?�7�q,��\��}�w�� Y��j�-l�R#*qK,�]��PH�i� �e}�?>�65�x3�<�N��L�"t�����,��K�K�Ŝ��6��}��/C�&�]I��?��Rw��֠qy�������vﰃ�����"؞˵��ևՊ!�M�N�E�d!k��7�&nF�"�x2s|�ҍ� �~l���~N53�0����ƥ�֓����s�N��o�Gۛ ���y��N�3ޮ����ğ�Ǎ� � ��}�:@Ѿ�M;ѐ	A;1_Z2*m7;޾V�0(;aI��", `�$j�/���%x��6���R�X��U��"�Lc��]P�࢈�틒+�f�{��8�^��6�[dd#�� ��V	O/�0ͻ��3�)��D���If�2]zQ�����oΤ��]�56���w���ͷ���0B�d5[�D8����4CL�5�g��s^�&�6��i���!I[���A(;i�~�F�C��i��9)�����ɬ��h��N��|f�����^ᜆ�>�W�CG.�y���أe��w�=<>���a�cz�f�n���n�1*ud��4Ҥ�b03VzۼAM/�&���T���� �5�UGq�����Md۷���S����#���x�g��VZ��C�^h�C�~�"g��hj2	�v&O��a:��nI�_�L�Gꔅ�66޹^�Xz�or�ZLK�YeH�9Qi�z�{�F,H��=��d&�%ɽ�+�'�ۍ��o��i6q6˺��#C<�]�@vlI��{�
��Ô�!�\�H���*����;�+N*����h�#��K��K�����o=x�#/8�� %6���C茓���ý���g�jEB�Z�b�ۅ�+Ef"���U=�*n�/�C�KqQ�@C��JwJ� ����j����>���WG�"�a����������ۆ��u��e��e4�Z�ċm��e�&G�'f8thb �#���M�A���+%��������o�f��6�e5N6��#�pI�x�y�WV���ƜĔ�W��^�u����Y2��^{����;�hZ�y�ʑ�����֥���p�L�7з��P	��L�+XC%�����ʈ�*cz��h �msg���Y����Ԭ�Y��|���Z0��D=B�| $"��#�h8���w�F�w���[��?(B���[�]"��q�Ce'.��c���;_G����\�̰�
���s ��;x����t�����W�[�Ѩ��<�!Z������ :LE������eXOh�%\�p�;
� ��bTe��mH�O-��I/t�<��'�_���GI/OVVW���/�Ī�BLJĢb�eI6�a̋�6ՙ����*y��D��D�(� �ee�#7�a�4�
�q��%,�
���5����Ri���� �S�fq�y�g	�1�.o�Bh��]�\�"l��ޒ�0`��PY�1�d�dM/�/�5�=�e�nP�Q;�>4dQ��o��k�\)�+,��(��j�0;�1�����xǼ�.�I5��k������]j��M����xɃR� z_4JL�~o�q����L�����L��8L��;�	g����r"������MSo+����s�Fvԟ��%K�p����z�����]��ꔽTds�� y�lcկ����1��������ǎ:e�U ـ7"�"Ľ��tW��l�v!�ÛF�����?��������_��\�����S�e�����li��t� �E�I��^���9�ղ����f#�/$������rxY�2��rܱ�n�Vᫍ4$���*��Z Bo`�a�kD�P���$�Ti�7��Y���j���oR�+N��L 
蟮��S\윤�|�_N��Ǎ+�����
�<��Q�_���G
�H�̂�Y;��uB�(�a�zS0&��G�gw�CwS�(�vP8O�.-���P��X�J��!��W^x#=��Y�h�5��l���I5���/FQ��
3m��ʷØ���oi�kK4�K����u�)������b�>sV�E�;�>��E��ka2o���n�'!g��0�l-}��gZ���<��!^�Â��v�n�<�B%�\ޤ�a�#��lO[`��$���D6��:�P�C�Kb.�����%�DH�;�O� ����h�:�O�>[9=�>��z���GY��7���x����ߌ�\�T��L��C[��_��E���f�:�C��S��Z[k�������Q�\א2��+��^ ��|~��Ok��`�T>�'�._w(��~���HJO��*B���c�/K�6���k�͇�HN�\������>��NK�LK=��~���Ék�t�	����!m����`3�4,U3����C_��S>�q�J�Lu�n�s�+
�Di�j�s����U�,���>��v(�J�Q�H����'�����v;�d�i�@6��hAS;1I�rq��t�T��:�4�	'W�Δ0����z�_���
*��S���l0�,��m��A�L���ՠ;�Ї����y0l�Ď8�/��ղr�
ѷ�i��#;"�q�����J���ց����sWg�&��da�-����]'��=���ag1ַg���������p�V2_Z����e
+Fc�l���'��a����@y��=�bT#����:K�#B��v2N�ɘ��{��&��.{��J�A��;��f��P��]���x{i�z���,i�>��j��F���;���L���F0LL9���n(t_)  1���ѹsN���Z� 4[�[`t�q�z�%��9�d(���#��$�x�,���q�i�\8���؟��큟�*���ŏ�-S�MP������&X�K�]"�?䣧�	(a���n�,� �<��0i.8%$�R�X.����Ҍ�w��H�\�5E���;�@O4����2�|Y�������m��\@��ӊ�*�0�_�r��M�l!¦Rh�i�vڵ��b=:�[r�2�0x�1Q���êX�N
�
=L�C��FØ6O�zφ�'g��5E�A5D!�%�b%�~�S��U���Jd����!�P\NO��M�Yl�B��U����M ��T �\Y%�Y��ن$4\G�^�`�\8[��^:�Eg�Z8��0ק�DK�;���B�K/;�=��b�ל��0�J�����s-ܵz\�*ڸuH`�V�k^:a]�[
ܾQ=�NM \��sh��E��H���ק�w0�Ž����}B�*���#�|E��^5�!��b��ڷ��z���P
($���T3�;��̖��.H_@����%#��Q�
wL�g��4+�+��j%�����',���VC,7q-�}�:	�*99L:��!P�|#�/2ٟԯl3g> �3B��UjXr�J}�6g�� ;Gg4���q!l�C��>eG�-�F+������a���꼃���~�T>�p.R�I[}�E֣JLS���j�{Z/۵���a���{�r����e�m�n��>�j���sJL�Ri6��Y-��?B���
�ǳ{����.z|��<U�+	�0j������ ��Ҹ�b�(53���̫���Ľs!�.��� �|�Dd{�0��v�^��B�҅��;�:����k�Ĉ�����LjӷP���^�(��nS(�8Xve��	���B�����|���]x��S�e 	���Fv��wx�ḁ�mlEݐ%W��n�l��sng�+�w�i�;������
(�t���)p0��,�ɢ��!`��)���l-�|o7x'?�>T���1�\%�J0��j��e)_�ߋ��� �j��s�N�e�+���s�e��j����7��~=�Τ��e��2R��. 2M(դz��C�V93���e(��Q��Y�hn��a魣O����lS
)ĄNw��V��[i18*��\3%4SR�3n�1�U�_���a0�wlG�b�����|�[��Dx�0banh��i?���1�3y�o@a��G�TK++�4H�yy�#�r�5�S+���w4�/3y��yZ֚��=n���7e5dj�xV�>�%^Ee��� l ڭ����?e��7H����|���dcy+�?u