XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��2!s���ӹ�E�F��3��p�k?�}V�"Ǎ�G�1GJ1D��7��:��;��T�� gz��󔂒�j;.��O�$�����-+�<Ҟ�� E�������W��m���<M�7������Y���ZL�\-\�D*���l���>��pCdנ�eF�z��s���1;����J���c�#����Q%�ZW}��r\u���c;&z?���3h�����v�0	�Dh���i�:���4�\eq���:AO�ґF�:��1���������0��֙�l�x>�w�ڂ��%STb�1U�n�k�G�t>6��eyx�Ne��m3E���˝�/_�����:p\v������S:�F�<�;#q�^�&��lL�3_f�I�R�Դ���)Pd/���A�"�4�Sg�E�-�8��n'��d�k�e���J�D��G�X�WصO�H�qU�Tbm�{'���,�21^G�����|��Qj�c��	��q�0k�X+�?���z4�p0���)� �`���U����}:r	Z#�!��G�꤇h0$;��w!��D��^�[o4SeE�y�UY�������u�N3£�����e"ɹ�xia�㉽�)V�dE�{�D����*�@����H.'����UE�t�2�����H�u�Z�B�U�VZuX��=�vx�F�u�Yx6��¤�1q��4#t8�����G��Hԅ��Jץ7��Bү���f�vJ�����^���E4����̹:�XlxVHYEB    88a6     d60<�*Ґ��nS��֭�B9VJ)��,|�:�jr7�"��+{�f\����	��5��#�� �(���ܢ��Smā��*��R��?��J��[�OI-r��x"$��	N�5P���R�3�Lx�*җ��&5�rD���kÂ_r�\�6�©��rȨR���p�;���,
x��@�E�45�$u@%������}g3b���]d�=��<�pء芁�B�`0pv�I��0���Z�=��v��)c{��G�Q��`G{f�1���
�"+R#-W��'��j�^/���NJ@Ѹ�O0#�j����'fd�0C� c!D��3�p���4g�]`� 1q؎�1}"s����MyY�]f7}�	<+ ǵ�m{bV�/�'�*��`���Xo~���<<T�-)ԯ�x&��?{U���DzT
�Z�J�K$�����;4�f^�ښ]5Z:+�D�H۹���^^`r}bR��NQ��u�AA6Y�Ѯrp���L��ᄻC@� �O�tpr�A�����;�?�F��^{�u\�������}���h�O������L���:�в�9H	-���ֽܜ�dr�͋����������;������0��åЍ����B�� *�������}��-们ǳj��;%�^NX�Gf��ԬS��璴�	�I��%)���3Ӱ3<Y�6��B<�y|v�}:���=�~�&X���������{eCYխ��6¹g�
ppvP�P�1�-���%BβW�Q&�/�ǧ��j����H��4���'��0�c�M��{+�Ӛ���6aKM#iw�&�"���d|�RzhO=� �	o�5����M2���+�w�}�X�|�����O��0,�K�za�0Q�(���S�+H�!��Ó������b�W6�K��fg��H*3��lm$�/�'q�v�P��Q76�Y�F�T��؝�fƚ��ݢ8��x=���%�����E($@}���Z��&�����;;f"Vz��f[JOGT~�d���њ�*��~ذ���!Ҍy(K���8T������+��/<��_�	�z+�v�ȵ��j8�ߕE�(n�[��KQAQ�F����2��]Y��G�~��s@Y��i�b&A�R���;�j&���&�mryҦf�n��GCK��� ^=*
X�8��u�?�z3S��0e��h�m��Ȳ��|��b��	��#OD�~?R4�+�p�&�g�Bt� q���"b�=;i���0$�֦*w��α��� ��Q�K����(����d�Ȕ������8��W�5���C�p�x�s,ג%��EC�⨸V�DiӦ��Eo^�״i|k M� Xȝ�h�oz��!�ۋ�-�ZuҤT��l-'T:uk܉�������Zb�d�\
����)k�{w�C�Aݓâ X�x.�k(����Ȁk�Ĭ��1/Jq��$I��E.����/�������I�l\ �!?�4Y����]�.�a��Aȥ�2�}�(���K���S����W�2J��HuƎR$��n��;�0�:��g�j1D�#|���y��wgLN���i*�L�$�Ⱦ�X@6�?N�� �hQ.�3�i��y&;��]�g����G@����Q��o�����3�'�m.m�b[q�5�ض!H;m�@S,-�_gq�m��%����C���-܇dL-�ҹ<\�Ы5s�X@
0G@��T_B �rg����#�q0-R� g�|����\���9X��4&�%��t�ki���q[z]���Ax1�a�DBء`�cR��Ƒ��=R8_F_�θv�Y#%�M �>R����lC�E�8�\Fw��[x@�0^^�Ǳ(��rOr�Sm�+j֯�3x�3���n��O��mK�����jgU/nwH�e��⥠p����	��'��M�(�o��YQ�r�Z����'�G����n����~���1zF����5"���W"���-�:����G���U]�:B&�ͱ�˜�Vw�b�pH�G�t�\_��g�C+��.n����_C$3�Vc%����I��
�v��6���5+��)ƒ.o5c���ѐ�j+���I�e�)�-n�QF���b����K��zw�ZR7�hK�IRUpo6�b���$mC���vRg��#�Xǳ���x���o���[����Oo0�{�H3�>�� ��K|p�aX�A_Ɗ�a�W�]�����:q\�<�!9�d$~b8���5H����f�����'��%0���;�2D�O��\g�p��9���]iUD�v��$-!{�VI�L���F�xc� ��eu�cnj߯,��DN�5�V�+�W�n������ %L�T?�EM�8��Jo�]��~A}m�~'�/�@@�����}�98�B����@ e�4���\����Ø��F�0:�wA��.u%\�-���cn��#`�)�kj�9/-�
��%H��nb��z�d�懯(	/HWiՀ�)��riaR���p芿��RszaN��d�kc��x\#�6+�@�Ӿ��pP鲒��ƢZr�\���] �����$+a�~s��/oX�<���L5;�߁��u��������zC�P!L+��H��:�U(d{���#�g�]���e�z�K�E�Q���\��S�&��7��C��l;vn`���a^QsZ����$����Uȝ�u}1"c@Nԙ �M�'�y¯{}�2�s�+C��90#xw/[]���e���zU�X#c��U�]=���(�� ��,�z&K��Dm@d�PC�V(���(�TjQ$����~?�fov��`�վV$:�+i0��u
ۿ\!0��sQ�'5��cj������~~�7�dv�1\+A��dEo^F.X$��@&"�{D�N�ڞ��m�H(���Ī��7B���JM�"�W�~{�C�ruu����B�>�[T2ok�l�潢��g49𔘊�X�)m$�
V#̤>�;D�/�+��j����jz?�|��Z1��;GrrA~{j'6����Ee��e��'�� A�9�.P�+�����B�~�u+Yis\i�R[�̮o��>����v��JD�_O�E����V�CT/mڱxf ��Y9�I$	$�Z+ r���,L�_)6�&V�ڱX���G��9���X���f�.�,�'�Bބk{���wp����|�,!�X(�(�S.�`�|��=�[#b�KB��>�oK�G�y<� 용3�i����r���j�E���ev����٨�<�'t�ѯL�O�/d����!�{{Ә�aO�1��+�p����El�I�8��J��2%7�#��r�P�'�0c]�eS̃�����m�ޯ���4p���g[���:����/E������*_1