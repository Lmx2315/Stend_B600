XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���@���|j��$�5��b�����G�,�:�I{�R�x�E�B�/h��\ꯎ{�?������G>q\+�j����f(�Р�jh�����x1�#m.�[�V�XT�7~�	�N�j�H��Q'���䣗f����͚��!+�.����$|�[�+�\�?�]�}�3!f#�לr`��8��v�[�k�D�0�.d�ݯVQN�M�?%M�9�קMnl
�D$[@a+���Dg_o��]P� �����~eO�I���Zl�-������5��j�M�s<-xCd�}uų)�3�?�#*��DZ�Fh�]����X�ӥ��{o�	W�f�4m��S+x0~��¹*��)�u��f�� �|�\�&���U�	��L�Þ�Z6�i}�W\ ���2�}=	�d�s�J��)��w�����5��hO��]V�`3�_A�!
�U	�A�$N+�ٹ�+�2\������ 8H7���>V��IGa5��u#������i!�-l���cS1DWyɾk�g�u)	3`_���8�Y,���J߂������?�7���L�_B4��8��,�u�ׄʽU3;S����م�el�顒07���7-(0�,���|��W��W:�t�s�B�gRC���k,����w/�X������Y�Na��o��9��E�kb�f���o�(��\ۏ���n��=��m���C�x�{�y���A�W�2|�V���%��ہ(:m+T/����x!�P���Z�ݤx���d-~�e����OJ�cXlxVHYEB    60e7     cd0~�H �b�xJǪ�pC���Y��9�j�t�+�Q��hwm��YGA�LN0�}v��Ř` ������;�4���Q�^�yDU !8�H�P@��^Ԏ�����5^+N�˴�v*W0r*��o�VNw�1��H��W�%�}H��,N�EZh�Թ�٨�J2xU���4�͑5��!|��A��
�`�����zM�Z���S�I��Ț�}��=pIr��g��֙gZ�|6�!E�]��c&����걒X�G��"@DI	>�>��z|�!��R㧷��%��o�����(��{XSAo��}�g��R���$�7^Ԫ���K3�w @���d���q}t�w6���O�Xf�Z���
.���9���j}��T�'t<�vG]�6���ǆ��sd�f`ߚ�*��מ8�P��w�'x)x&N׵(u��M�%���	g�e.���ڰa�U��s�F�$�7N�;�����W�'~�{
�E���$	�LC��چ9|\�#S���!+�4G��[ZÕ1�Ҋ Q�,�4>gnO[�Н��jka��2��p������u��V.J����y�4f�F�C�|��09��F\����]�]����I/@���ߵ�=�LJ+��n���㊒�x���E���C�.���GC~�Jf��Ħ�v�p�m���9����z`�.\�����[��>S�{2�`b�H���^
�W_ �M���M���KF:�r�Z��Fn��[��Q�)�癘gC0غ�⊖/[ee�m�\�)<����k�DS7#M����r��j�^�8�z�Fg��������Q��b��,��bLO�Z���i��c*��Dq��I�����o\YX��[��~��K�J/��玔�eg5%�M)�G� FS|J1'�=UDh�>~uB+�V��{�jGŪ�&���~���}�u���������U�V��O�VH��QȼKu�}c`^�/�P����]�Qf����y�H�+�\`5�;�'�vX+\QU�
oQ�UdU���Ś��p�5xsJ|0�u/�=GD�@���6L����G��`!g_�Y�U��g*�](Jge `�U�Y+ ���iƨ�� +�(MZ�G`�K!���.ܨR����B��ƃ�jeNߙ�`�W��I�B�n����S���0����	�L���e�6Y�;��|Ƭ��M ������Ya�S����^p�r��!P��MT%+��Sm V�W�B���B��M�e��`�}M�PT��V��$��������w��:����w���Ʈ���`٬t�ڬ�Rg�:��p���>�
�K>D_Zp�<(~��n��UM��bqp�s�j�>
\�^:�RX`�;��δ�>�
T4�C6��_*Z�s�Ѽ��^O��R��WC�D�l���y��O��9�ѯ�υ)Q�أ��M�L�;�T�(��q	W:�h+�E�#��-���`�F�ƅ��L��(��P6����n��A�ӎuᜰ7��lTZv��j �d4ݰx��j�����e��xI� ?�U'���$�K��!)�Z�y��GS���̙�ʐ�-ރ:�S��m	M��9�'���_X*�(֗����������6ՠ&K�$I����׭U2=�A+�>U%�gEWҿ��;~�;�����^���,�U��L�$�I�[�ϲ���e�����5F.�X�%�+�jX�	5e���N��9����P! ���0��@�O�|݆��n蘩��	cs���#��WJ�[�rE��Y��k�Ö�\�{���y�h���fƥ���x�I��Ԋ�8ld��C)�ZAEV+ؒ"�w�Q��r��� y���xd�s>_���(�4�j�'���Eshĩ9B�
F�J^ DX�9�-�M|y&��;PX��g�V~h��9U��B�S��A&���KO
��Ñ ����R(t6��n�2�K�i�RgT�C��,(Β�^�&��A�a��,g��3jx��1M	5O�}�d�3�Q���l�."��l/��6�W����(�]���tx�/�wb�ۼ(�`�5�p��SS����:�������Β��9�蘽H�-���(�I�Zi�g��Z���jq.��D�oo.N.G}�ўu�v�Nv9�Ts��=Eb׼2�A�g~�Z�>��I,�$K�W��p4�kI>����������Փta��t�_��N�++������M�cbm��*�k�	���2�#��?�uy|%��Z�������4�+ePR�K?����o5���Jߜ�0�p�lt�&��D�}����
��%�K��������x���渰��){�uIe9���
��`�J}){hom���-�ހxK����*�|��VW�-��l�M�G%����S�tX��l�I/�:헁�3/�?���'�1�Gk[x�pcJ��X��Ct]l�[���0�1����G9h_D�ʏ����z���J���F���V �!�u4Uo��ϯ���E�@�X�u�P���}d���u~�/����Y���JC���8_���2,-_G�k�߲ͯ���f|Ȏz[l��x��U���@qe���2ut��
��(�����ð�"!�_����nw��t�2�e��怭ݑ�����$��J&`��z��.�x� ��GQO��k�qpv�zl_�r2ʉvh�����f^1gO�k1MQ֎[������_Zh�x�
8��kH����8�:*��P���o�W�x~U0���T�2v�<")�1�b����ͤ4G�>Pț���ʾ۪��~J����R_�ի���̠X��H^s��j�&�D{s	�hB��w�4��� �|]��c���D�<MvO���X;h��8e�2�N9s0;�t,��y2P)��H#�VPQ&[+/1�B����&|��2<P��T���5�h��%�HwN �ͨ�(>g�}��_��g�r"���d�]7c�����q�M;�2}���@ZYb�
����Mo2ͮ'/�Ҡ�\ϗ�S��7;����y٭̣T!���ZEX&p,]��+����K���hyS�O�
f��o@�*(�s!�<�0˸�yF2R�ͺ	�2s��"�/�#-�(
a��A�����GL�X�mn!֮�'s�� d�j\���އ��th�!��$ݔS�6��ؙ�̏/�pb��u��P^��J�v�:��T���l�^�̕�n��F6�7��