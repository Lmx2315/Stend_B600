XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��]2�k���I/FM��x#����E�.9���C>d]�����,���V�b������QE�9�@	@�-�D��u0�Az�;�3�V�m&�/���%
˭=�=�_����~���rR�4cg��3.�H"����	Nv���m`u<�`���Y�i惐3<�	��ӫ�Ab�g��4�E6>ȍ�!׼A)&�� ��iȕ�d�	�)�{ �c�c�,$���N�_ VO�1rc1F��?m�]�~2�4Z::G��fWUo1:7�K�d��c�J�v��?
?iᚽ��A�S�䩏%�~�ϡA�Ts��I�T�yJ=ߗ(�y�RvӮ6�o�	_ �
U[C��v@�ǖ^8ǦQ���B}���2��	ƦFX0@}"��5Mw��|���Vf���"�Z=����]g�
!�ս14]7���설�HQ$S	��0`h�GF%c>��wv)�l1I�F�vH;Z��6L�J|jW�W�:�
����|���_S�u�+�h���Ґy7ˋ�#@�tKA-����V\A�0Ć�����/:�ج���Z�����]��M�ۉo:�.#����7�"�/� f7)$H��V�ꭗ����/��˺�����.�n��\`Ʋ�׬!9^$(��3U�<����u��)B������NF���]�퟇w�qO���&����h��q�b�����\<'|ވD���Ϻ&�Y3���e�ſ�Mwa��9��{���RI�vyD�_�s�� �^�ƀ�;$P1wfr�v�+Z����XlxVHYEB    41b6     c40�?m���η`������Z���a�/
et��i��āϑ9��ܷ��IJ<��I4��5������V�Wf	�����H�dwT����5���,�a!@G|C'\��U��?��E@�UH���4'�f4l�ݪiT��5C�A]w
����]��9ܶ=V�T�0�mg�˄s����b��q������A�@.����y!����O����ɒ2�\�W�d.�_D�������O�ė%�\	�L$��i^�X)#�ľ"7����}�L����asЎ��הZM��э^5e��o�F[{�!G��	�M6?K�P�&rV���j�F(�t��]�þ�A;��ޱR�|E]��p\i��ɤd���:m#�E�\���~vLK-ɑ�9�'Ȧt
�o�i1n#�����hy�,u��9�6�4�����1���Oh2T����nbe�R���9�4��5C
��R�u�w/�[ZC��P24A�9��
�;�Rx��P ������J�g.� M�& ����42s�Fg��������y�nv{]�g���-��p$�BW��Bsy�
g|]w�b�	L19x	������Q����"<�(U���g���+�7</�W?-Ĭ�r�J������
��z�#�L~?e�/�b�9k�L�������ظ{3\��⍽C��Y�7&�  e �%�K��N�I}�ע}U������P�k~3!���g;��]��

�qz�<8�P-&I}MHSҚy�A���G	)����s�F9+מSI$��A�k�,��j}��?,wS*8��q������;:׈�[sPj��j��(~��ب��ӣܼ��4�� T�X)�>�4���B�ݕ�C��C��u��	;d*��cTZ3 ���q?}�E��8��;~�a'������Ӣ0��L��_�wX,3�H�7799BX�m��+ v���BG尰���ߑ��M-��R%ҙv�(_ހ"�YR`UP��h��+���D�x�>��e���0���ܫȷ��ݒ~H4Ioo�@�(;�E~ԋ�s��6b����;s��%2�Q�����9苑e2�Gd�Bm�_�D�3�4B�M8T�w�ZA#Va�907������ܜ6��ē,��K�OO������r���t#!J�7�!N�'IȾ�];���U�gU����`�������#�	3k) V��T�KV�Hq�8�fe�W(�0!�Ҧ�`��8�i��Y�@�:�~/�KB�{�7@�-����C��^���f�����p䜩d� �[�â;�K�>��)�����z�+r��q<�#r�A�R��z��BHkƘĒ�i[�	�#���`���F���&$��Md-"n�#f���Zx��x��7s�`���}��#'�G�h��B�؝���Ne������.�̷���&��õ3��C��k�cKЀ��ߚ��v=�F�dzg{c�g�����T�� Y�(l�s��!��] �[�jF�f�íʣ�OS��r-�����f j�{7�40�	�f�~���lZ"l5�*��b�u#q��r9�x\��nwґ�:�hౄ��]̠������fvn��u��J�'�K�yO���Qf��oɼ�<�B^��X���)�T�eԿ4;������@�� #c�6�;�k��E��k�G��aB6��r�r%���ϭL��,G�V�p��V�a�ª����%�[���"v5(�m�f�v
��&���4dD���;P�H���j8���������Y��L�~x����[r��i8Z>�D�@J�H	8�T���<<7eސ�		7���#�x�T�ig���!'�}]?-�/AQ*�I�Fd;T����Э����xJ��y�2�Q���,%Y���?y@� ���ͨ�٧�����1�U����J��S�5��4�e���{�]ʸ�~|�U�M��j8�����z�]�B�}�lj6`m����	�S�V�/)P�10���<i���a�����
�[b��2� 'J��LI\��-��h�h!�� T<��2����E}�;>���b�/!l����N+X!x�ZӤ]�Z�5�יcfB���IH$*)�E�����	�u2h�bK�X�΢.��1!j�i��~xk1S���@Y-~	�$�׃���2���V�������<���J_�� qiZ���H�~��M����@�.jsoV�D��v���5~S�-�1�K�����)������lx���輻O�;�[�D��VX��!��~�!\���-��;VU<�h������s�GϨkǵ瘌�������j	��	Jv��_6�F ���؏�K��+��F�D[S��IZ��8�֕azX�`3\࣋bV<0�Q�[C�~Ƃ|r��~�mw�T�ܼ`���zJ@�ؿe�L��ϒ��*�;�¦ۙ��k��݇�gN�x ��U��7$�"�������-�s�oH�7g�?��pEM#���(�oe�n4@w���VM����J��9���J>��R�Q��*=sf�G�O_�/X�������[���L��CE�N�B�p��H�/f˙n�qڗ�U�@j��8!�e�?ga�M��;��҈�6�8���
4�ԃ9�`R�2۽H����|�z��+��,�C�^Cy�����Jk�0!*��*JRN�d��^�I�?%��d�h�۵l2u��Q�����"�E��ㄉ�׌��">h]d7�}]S=e��'cgd<���T�i �Z��j�\��M���9Dr_��a�4�1p!���e�e4 92��}������m`mX%�>��W�[3A@:	NgvT#h��L]��-�M�5���s�o��Ս� �
�S <�EK��GH!-ܛ�����˰mЉ���}-�>K��3/�<Gc6VA1��cW;G�j.�S+p�b� ��it�T֡qb?FM���aMv0*l���Yه�|i���0:��j�Wj�Π0�@�k?f&��f3.]��źbY�huI�LN�ZV|-���~�L ��5���3D4H[-�G�Sy�r>��;]]fuX����g$�2�(��8����e��e}