XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��S��������7�#J�����8k�����]C�'
�x�'*�A��=�Μ��%yR�S�:k���h�/��4�� �q���RsR�Z97��S��s���r�&cz�AH �* a�H��wT{�D{�y�J�GL���l� }_�Rf[���&�&�Q��Ъ%���kJ���g&
[>���?�q<9�/���0�k}�3���\�(g��ӞM#�� J����'����)u1n����?�F���+/��y���w�eT�6���+Y�I$슃T�Ӧ6��d���!9]Q@���s�����°dS�XV:��eL�cZ����{�)��?�e��(�ͱk{�U��1ʝ�ww�
���[����r�>����02ރǀٍ���T��E���/�h��ʳ4�W��a�xB���������Dm��$�M�BJ�T�h�f5Ζ��z���g]�b�H�=�)RPI�T�(5I�]����4 ��{���?�S�@rB��j��;�YU��~�Y8~���GS��c-� �����G>d%��dJ��V�XC�*|����S9Fשׁ%x��j�.�$I�De���JAn�OR���a�	4X�a|7����/�m����W�`�7��xH^��$Ϥ��/6ד7�%C��,�c�T������G��/�����h
1�_AϹ��徵|%�¡8$�[��F�Y�h�K���TΔ�>g\#�\rh2,�\��*���s�!|��@��XlxVHYEB    165c     4005�UX�K$�b;�G��d��V0F�z�2|�y�E��T3d'g���]0,1N�p�5_�g^\$7�d%��R�)k���R�:!6e	9}�տ5�ue�1B���ö�"��IJxm~|����Xd
����\����o�m8mJva�@���!'c�|�//����/�	�g��1d7����C�;K5��������He�/� p�� x���)@P4V��-/���d��H97�O^r��G��T�-vy�F~ڱ�r=tL{�uG�?IB�GZ+��������%`������u�i �
��(�/I����6��-s��iV��Gh�\��N_N@Ү�����9��N�{�� {�.��F]�L��<�a^* \��*��Ϭ+�,c��,ۺ�)��(�pѩ�z�J ��\LLE_j�5Ne���sR��{�;�f5"w�Nƥ7ܚ�_���*c��4��V�m�'��[),���T��s�+�X�ή��oͮ���y����ၬ��������GgM�v�)�g��/�ڐ��g�t�����n�9���(� 0j�r�g�q��`��sA&�sM����5Г�=�zvA�P��]�@vZp�$r�<{;�oƭ����Cr,�-��ڍ����G�y|��(��Pp��V��/W2���y��4��Z��"�-��x�};�`����y��l����b���,}�a�SbW�!��u��*�9<�R��U��ވ����O
=
��9���}~JÒ�%�k��+�@�",t,�����Ƅ���g|ލ�S*�.���>�ކs��,l�r�
�7�����STT(��b��(Թ��pK���թSGh�
�[����Lt7Z�zlTf�ݹ4�`�֣�������� 5��7<���e��$NT�[������؟���j���3�B���zf?o^�T�!(��R���yI2��Yw5y]�{5暞:KBZ"��$��ò_r}V|�%qk��e���?����8�Tm��3g��4}�7`