XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��>�S��E"�����Y�>�l6�Y/���=�2
U�_ܸ�g��l�d�A��_�Z�Ή�̝�ͧ��x�rs�K��o�UIA�7U���򶌑��*��	��RU�V��p��4�=�hoR֕q��K�@�����:~��F�`I���_X�.�at��y�w����{�0���ڢ�_��I���2�vY��Xq[��@K�Y���d�6�w��ESVC��M��s
K��6�(F���-Þ�D��MnlM{C�Y�Ϟ
��h	6?i���m�i�Ch�p�_Ǣ:lq����H3>G��0W:�j��+vٕǀv� rw@FE�Ԩd��?hE�S�i��T�|x˖/&�,�/Png���y_�ϑ��jL{�nH��������Vq��_�����f�N�H.���7���"�n��1��i܎�A�Ahe,�Yw.(�+�o�符�0� T�j]���:��D4 ������0�Bq���_M�'C�����T�튺���R��)Y%����k��뚻OD"����_�q/���Agsڤ�R����3��THJ��-4���P��WٚؿS\����c"��2Cl����},�sD[��*@��E[��_����E��*���dS�r�_�ǲ�u�$� ڞl�=���?�5�B|3d�\G�D�*a���(wC�iA�F�!݆O��W,cL��Ɏ����sA�·�qFj�Cu��cN@��b�i�8"H�x�)i#�*���z�y��I�~_c��`,��q��f�XlxVHYEB    a6c0    1b00RC�17ع8�u_&�@C8��Q���b�&Nz����E.TQ�pC5j�Q	�G��x��%�;Bn$w�p�T�ݿ��5���}��J0/�|�ya;GI�?�iEKk��7��J�� 
1�� ��4yY���0_
%R-�B<���t�&!D�!���E�h�S;x�����	��H�X��x`�(]��������L����e�cY�x�d����*&��g��ˉ��˗K:N_*�c�q����P�������6��/Y�7xgb����:3��\&�v����s�=���R}�U�%���M�:i�1ݘ�����,�����eRh21S�ɳ.`�z���=G��C��`�ᡠ��H���a|�xW4"9��˿Ik�
8Z��x$^�v�g7��z-�nI�s1�ы����S�z���|' �9�i|����N��X\�<�㥥9ڥ;�6nX��5����9ш!ojN@��$�sZ^�3G�lӛM��SP)�ք�0�ţЎ�߹H�U���s?�B��Z�d�SX������Fm��O�=(t<Y�;&-\�:��*7��bN�#;�@�H�[J�;M7&�)i<!������qG����%@|W�bx�&N`� �$9 ��h�	's�5H䒿d~vS7M��<�6	�����/����eQ�$9��9��ط�̵�`׷��|@lWz�Ѽx��>�pbg�iX���)&�B���Ω�,�3�Ear_�YGV��IQ��9��z��0����%~�0��̉Օ>�Hi�יA�ƈ���%kA3Gp�j' �)�#�i��������c �`�eN���ƪ�/*�"�*�\J�k �A���+�L�}F\h�y�	�1�7�S�I��P����f�������k����%W]���s˿6 ��~�	X��}�Qom_5n�V+���o;����ʹ��~��G��E�Ax�V�Ҍ:��v&�i}�I��w���{�&�'�����ٶ@\c�Y��ߛK<8�M߄���_�W"̸�ڑ��V�U��c�&
�]��Q��D�(��e���5"�D}�g���]u%{���Y�N�%3���I� �|��x�Cc�sK�""�����%yjw[p�Cz�L3��G8L���$H��p��dј9�3������&C�)	��B?��{\�� ��Ƌ"�m,A��J��D���l���r�R��0�$�[K���%�j�)AF�ao����3�Q?�NH��LH>5~�)��6�K�Z*V|Tܗ��Cr!i>f��(ղ�Wu�t�~��s����1�&cɌ�L��k7	*÷%�\�wۧ��z��ٜ �b$���s�9[�V��`��9�W|у@�1!���.�T�q]�|-Z�xG�I��������
�=�O�+X >��R .K��K�~�	N��>��Y��O=��Iu0�N
��2�7���n(��]�*kZ�F@;$E��Uҁ�t���]!&�<iw���C��w��k6�l	���_���և#(��d\P29D������R>ɧ�����<p���Z7B���=|Rö�.�x�L��#*6�������_�������s#�U����:��3n�?��f�~�C����Ci̸蔺,��_�/�T%��ٸ_Ք�7�Ps;:���6��r��ّ��HE=�b��ט�D��d�{bO2�0���^�e)0�qkUC�
��ڦ��Ԗ����R�	Ʈ�
�e@�4���ҏ;׃��?~[�K�YQ+��I�.������R/��%�n�-�t8��%t�:R\IZ9��5��^?���j��`نY_���H,;���G��엹��4��yh�0�+�#�M1���K�����`r�]����0?q"�]�����N�0x�\��1x���mЄ�\ Y��
��/�׳�iI`L�50W������P���g��I@�Ҏ;�6�K���q�-$��#nf��wp��V�ɿE=;A-�Uю���������ݙQBm��de"?�{���Fȋ�7j�#��^�+]Ξ�S�_�~5i��������K��BYo���x꒸Z�V��%3z�~M��0~��i��ˎ���Z��������}�М���뻙�7S`����R�Y���p}�-	CS`��j_�g\r�,�^%�ñ7)Z��l6���$�j�m1[�	�D�9�������	�zj:���/@¥%,�D`����vEL��oh`�_A;�ڬ�*'�+�V�1۰��P�d`��Y-�����՘�p~7������h�y̎$��e
��o|.&���l���HJyV����a;���} ���k��)+X���e���� K^	\�A�����^�@�����[����d*=S����9���=<���򢓛F�b�A����8L����/�=Qˍ�]��t��Y�R�陗{�ק<�'86ӄ< �Iq��Ȳz�!��W��5f�1������H p�6�Sm���;�>�1ן ��lLMxx�����+m>3T.J��o�H7��s��^S�,SpҎ�3"`��Q�(���i�:���ګ�l��l.\�X.�y�7k���h����J�.���_���K*2Km�i���\x��t����}�.��*��x�\yL��g�Ñ��^[Ai��o3Q�����E�������ƒ34j2g�P	&'��"�At�ǳlSƱ�-p���]B�M��<�7��jqB���p@��/�U
'��gu3Um�b���Ga�Y��)gk�|�#�l�ҍ0�(=`�`�,�&ѫ
�B����` �[�W�`�$��QJ��"+a�Q�?qZ�訶X`�\	*l;��W:�p}��ڋ��j
�
]��� �	��X��߈b��\&B_��~v�B.��a@9h��~��yEF���H����'��E}޲�h`��ԓ"%Z<�=��g=0p�n�+�&{e� ���7�ܵϕ]�@=�P��M~]��&��&��9��XX�&�����N�t��E�����i�"��( �S�!�4x�̌9�Tu���C����G��	��X����I^!`��Ƙ����S�}��j_'��؈���rn�
��\�������ĝ��d�<��/����/��g�<ի��7e���G�dL�t�u��m�ẟE�}�a�"'Z�cI���h>��5l�n)��5w�����\��l�Z1��o�c�eAE�vM��9	�� �K\�l���=�㾰Q�u��<�FP1�6< v�剝���Hc����m�$���m�U�h��*��;�]��&s|Lm��M�`<��j��C�l��x��}����k#2�k��f��E���&yv 49�~G4�H� óh�q8� �J��*�L���k����q;�&i&�^BY��F�B�D�g�2G�)�G�-�e!n���}��W���,��}�sKՂ��Ż	�q/n��&���΋�&PTv��k{ab.e쑗������ā?��p-^Q�-F�bt���Z�h��0�fa&?bL�X�@x�(��a���@��\`���A

���z�J� �E4�NǓ:ǮV�����1`�� *�6
]��7��kX���J����� ȹ��1���s����ct��#���6W&yY��p%���9�dQ�� ��m�#���~_+�q�����+Q���n��@@���c��RSo#Q���yq�]�V��f��6*dO�l>�*?��Ӽ�Ti٪q�;L.��YP�T�g���g2? �o��0���$�HG[f��@%�����LR2*B� �T���L����N-
�|��wh%��$E�����? �P���Uʀm:����*��8b�,,:'azM�S�z��|�х�N5�����Wb�8�`ٓ\�e�Q�G����p��;�55�ߎ��c��װ�F��$��Rܯ`I-Ռ�ʿvJ�'[��@�*8��kz(�{�u�>����F���[��s[��X��KG�o��H�����ft�p~, �.V��{�I�ݒ��[m�O��%d��JD��i�H�<�ձc��t�Z��o����Q�s�l�PgB;1���7#2�(h�K�k/:X�O���	>�t�qq:DM�v܁I��@�c�~�S�$r�~,<�g��Oj��;��k��=��F���E���{��8�/d�FU��6c{���1ଗ�:>�	zJ8��[k�y�3*�@W��Ah��1�˪bC&���:�}k+7���ږ�5kF��l�T��D��G*+�^�MB��,ȕ�� 	]4�.e�h���ڨ�J4j�n�&��X���v��B�]m>Y��I+��ˉ���;���̅��>��L�8t�zِ\)O��j��@�S���1��P��8+���`C�m�+d!�:�}įyf���o�Qx�L�>��GqC�.����$��;%��C���-��LpL4A�����z`r�UD�6�����}=��EvG��5�ك�t}�u�khA��Q�6�&�ڐ�+}��g��s��]�,P�Qnځix��8R
����q��T�f@A��%;DS�|ܟJaE숖��	����W�-l���@H�k0	<�[�Zb �v1O�k,d�����3r�"7B��r��Єh	���ME�O�<�~���dO>��i}�	S^aoK��P�^�?b��V1j;�t<~�w*8oQ��w���r��^�Fj�r���6�ϔ�a�A����=�d����z	S8C�����+����=n���Dͽ_k�CUF�x��8�4�z+�S�]�Xf��2(�\0Ͱ��@(�-yѵN ��jƀ��<��J]K�����՚fO�S8��c����܇�D���F��2m��<����}�������7M�A ��¨��"����}��]eC��,��T��Zv�)&p�\� e3�C�#1'6��r�n+���c���K�~=Re��$�B�Po�h�|�c��kU�E������i�΋�Z.ߋ�~Je��#}
��,0��a���s�X��y��ujp/�����t?��ޙ�־"ſ�%'�M��M���̹�L�'V�w�[zo�1Nl���ŃA	����ō9������s�.�#c����:vɜ��v&�}n�)�H�ˎA;u�Ġ.��v��gU�/I7WHT�\��'��q"hR��s��ڴ����q���Es`��1D1�dt���"I���Zi\_�	�2���h䐓�aQ�S=��0�C��}��E\
�o D���o4�%��7N��Wu�x�9�#���:�8~�_�Jk��Z�b��b�����{�n���̲�t-��Ct�^Zr�hGq*�I��[��;��j,"��j�%�x��nn.a���eh_�?{�-=�ZURxr}�D�Ľ��d�gD��xM�_'��~�n�M�P����k��}����i4���9��T�L����z6"�?B�2F6R���?٠�.Y�%�>c�}�e��:wzo9����W���p�綄��V��}T��Ӫ�m�<���_.+����������#�mX���T�����QBx�����*"�M|s�.���0�cٴ��qٕ��ˡ�I������r�W0xi�ٌ��5�Ǌz6�V��5�/V�ޗ��N����_;}��Y}R��S���&!
v�ް��r�s��U~;�h��w���J8���"R��)��=����*d���X/�b�Ň���l���;��~��숺�sN���힦=�����E��'�p��S�>�׆�8�rvォ�J��� �K�f���,"�fFuJ�xny���jiW�^Q��aS�����}h� H�5��>�9����@l���`��W��R�/���$lټ^�A����4��[Aܴ3d��|�v<����e�~��6���r��}�K<��v6,�5����O���L���W����h����"��+��h�i�Vٽа���/�W��_���4&5HM/��^��w(��"!�Ĳ���4ċ��ڱs�Է���q�,Y��V ���v��W���4o4\Q
�l+��g��Ɇя�Xg�V��s�X�4�=\�_8��",��x�[o���]`������N��S1<5pv�����:X�b/t�D��W�c̤����R�N��ě��L�U*�*���;r{��+p�Ǆ##щ<�`������K�&����f��S�ћ�`�2�h��j���޼Z�ͬ�,�Ϲ	�QVI���T�H�"��ʶӹ��[M����C3��{�B���-�A����+:]h��#�)��*�A:R��fa�9�LB4f�2�,�J�DL��0|��S$���������Pi �
/�\l�p�l����R���N��ET+�w�����_��
���TK��v/��H5*���Q�`.Y���,\�ji��_�F�����&���+7�)�G�9�)%�D��y(�һ�¤���3i���Xނ[���H���lR��T�M�x���o�YI.Oo�p�\[�d���#���O���d��M��3�ٽD�15��<�����,�?@g����uf|���Tp�"�%�-򤃂��؛r�	s�U_�2��{�8�e�T�3j�Brh�n�fO22g�j!���}��Q�7��7����!���t��v����˿���p�r'B^9�Q:�˩[�k���c֢���5�Cp4����3"8�Xh��ʷ�>Y��q�q��j$2L�!�T7�*���1��0\��E����?��lT�Eg�b �C8�m�s���4D$�@��0���{����S��*�z~P �B��pD�� ��j�g1�N3B��M�(+�(P�`;�n�ު�Kݭ�