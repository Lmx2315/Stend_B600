XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���kr�&�{*�I��;k0��2����k��*��2��~���WW��DzS������a�A��K����W����Ja�8��k��;3/�mX	���p��/#�U�ڹ�/���{t�4!V�sy��}A�È{�d���r��P�W�2��	;]��n	>���>��&��wߎ뎈 �P`�����H�,[����#@��@�1�Q}�_�Ҕ��!��p���쨧�='��a���kꖈ��AX���jd�/�=�94�]���u.����{E����Q\5xΕ<����+����L/���󢡌.|�6!LX�����Y��~:C�C��z���2�PBy�a�g�!�u�П �a~��3}S�ΟMŒ��ѝE��{;���p)Zz�"��������2��i��P�Ú`�m�f�a<��@&s{ �	�bu�v�Q����K�HԚa�jQp�(��m�6�����J�&F����\K�'w���Gy�oT"$��,ePI�S�Nm�����*�e���t��"�&�ћIێ>��<ܵSz����%\Yo��F���w,I��J�X�I�q�f����F�T�����3�R#$!��+vA"��[b�mJCpBCꋡ�2��(�pVUnJ|<<�ip�	PBK7S�p>B)a-�z�g�#����7�˧-�[��^�q�xK{?���J�͝��;�Ja��fQ�a�}Cb��,j0��I1 ���`n�yV�=���
x�XlxVHYEB    17a1     680�5��Cj*%7c1���.�q����д�j%���< �y������K��Ʒ�b��jr��P�m�Uq��[�d� ��$�dK�X�F㿍�켹�u�:4М�jjV���D<��?����8��5�MI�G�'���g[������P��¦�{��A�3��K���c�9�gO]͑��R�c-�p@|��Z�']�ͼ��`J:i.�����y�߼�`f@�:5��1�I�xy|�c΄�F�w2�[�xB*gr��9 x�57�в�{���h<luY�k?��/�4{o�f,�l\��<�AaÊLH'�`��
�3ƹ��Eq��'t��'lh�8���>Qu"��*��$��f?�d�j��;N˯z��F$�u��ծU� ���R�Np+=��."�/�����Ư��q��(��}��x�J9����w����C9{����`�vY�,uX���.�8��X�Y�Ь�	���"(_�VLx�����Mn��������j�7��It.|��'1��L7�L� t��d�x�_�o��q|V�1��&OVڍ"��T�o�Y�@�Ҳݫ-s�Q�J'㴌�HFF]V�� FX��Jv�-���������jK��NB率Y�#���U�N�6,�4w[do'�'��͍7����'���܊/��(�;���R�9�{��1O O�W�Z�߅��~��h�VV�(	��R��E �[$��B���)�+p�o�{��yﯡ�'{�@�\/�n����c�,��лצ!oG��	
�E�Lh�q.EKX�G�AVC���BՄ� E����8��Q7wX?'吞�q��z���7-�V�����J*L�	�9�&Ϣ��F̚��PY�uPB��|𭋣/"8H�+g奓������U�pηdP% ��oS������ӧy��S}*(~�n^%o����	ji�j_�GN/�.a�L��+�̳�0�E�)��N~�y�z�Ʀ�)^c�:քi~�Fɏ�T�C-��dP�Dw�2���'n����p=��g�*:�o
E�A�v,���"v���y�g���NU��=s��::V�XwW����ǅt��E,�W��3�B���j��Q�-2L��6���X��P�֢7+)?�^�  &�I�4E�<0�,i��]S�P{W�a�@+)Z�	�l��S���Y��8ʲ��f	�+��N f��t�l��D����*�����_���yJ.s�J+(XN��7�J�\E6��<�y�'�K���՞d��[>]N9����`Ԧ��v�AQ$��!�F�v����z}2|��ct�������f�LO��(&��^�+"�85�H�S5g�-������ޫJ:n�G������c,��/v~h��d�G\��3����>h40�a�,@ �V�J�����r�z"�1h�Y�=;��s�S���J�M��`)��� �Qp׎�p����G�,�'��{��ߚ�"�MK�N�?]�X��������PI<{�C�F��0t�B���K����G��W^� Fhe-�D`U�1rP�lT�O��_W�U�)�O��y�N32A�|f�j�p>�'�^�{?+�2kB$)q{_D̵[׫!
�x�n�[8�~����`M�^{)޼#/��u�[�Z