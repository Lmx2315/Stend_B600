XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��#�$%Kʪ-���w���pm�[��V6m�
?�;��
�v�\f���,�������IH�j"I�.�l7��[?�
��OTT@a�@�l̉��K�+(�u�9�]&���|ت&p�7�����ψ��<��Y�<L�Nh��X�ɸ�4�}������H�ةx���~�%����P��!.t����%>k�'�g�2����85iG�4��^��I��p�hF�>ڊ�x�`D"�Fȋ��Eh'��{r�ϊ��|�G3�<c/oq-L 68t9�e�A�dx��s ï�B��V�I��MUt�7��@�Uĝd�p��$c�@������)�!E[C����#���6��F��;����E˻�Y-��	�2��.�oA�Q��Sm�z	R����.����2F��U�v�� ���v$��*U(f�v���Q��k��sη������UFG:�xxо����Z� �zu����"��Ȇ���Vs��JG�μ�*�vߴs��	ݓ�$���1�x
?�̪Em�"���NL�G�\K'��U�&[U��t�ZI/<�����n���{��L1I�f��/v�d���ސ�8�r������-�,A���ؖaXtk�;i׋fߜ��@��
}[GR���^hGbE�eT�7uRK4�!�t֫qf����9�IM�x�ie�p��l/�K��������p�=c��N�6�Q���eL.,1~`p�$sƀ�����O.�'*.�<�룄o����XlxVHYEB    fa00    1a50�,_��ӹ!����=���z{/�?$����i�!�㓎��O?���X���t���C?�S�F;��AbT��V���$kI����BF�$�G���k�/=��+)�#��iϵ��w���$~��{�X�����#I �r�U��{ϴ�]Das.�)�QRIJ�6��+�N)~T��t{�MK���+��0A�y%��̙1�Mi��1�D�L��#�8)C����ܭm��س�-d�N��Oy� ���6mhjah���\���/*�����S��,�f��!��(o�.T�[�}>0{>�h�鷇H^�~��T$g+�N�!�8n�f�L�,�LI��<�%6�Z;�ь��Aj����Ny���d��U��BE|=R���L�m�'Z,"$�k�
Ѳ�#Q%(�p��ּE�"��z{h�h='T����������u"�L��	L7��y�?�{�#���RR
Y�3o��"Qj�3�q���8�F���#���V��p�������W{�p�����%i�:�-o,�G<P�����n]F��`�L���/Q�I]�2a�xʤА8`Ǫd0^�jmi^2�^����m�T�@(r�9�g\H��%��Ǥ5���m���t%��yz���$T^3�����\;��3��&Tr7zٳo�T�w­H�mىpO7n�4Dǃ�3�����C�&?A|�8�V��C7ig��)�4���/��"@;�ټ��]||4	_�CvErJO����ݰcA��G�)�s��DTuc�gE��S>��֡*&��8�,M��>Oֻ�����w4��~�&�gs�?2$�֔��L��<eQ���b4���,��1��|�t���e�2�+:�F%�D#*�8��12��M���إ<o1kbې��!�Pb�er���jwt�9G�����b/a�S-����A��0] ��?=0����C���`�7d�U�{?�┊�3�v@� ê���C(_eWӒ��i���R�"�z����q�n>t��N��d���5���W�av�"`�$�K��F�>�E��e��9����5t"E>j۹����8��cz&�u����bAoڑ���;瑇ľ1"�?}y����ťf���7����?���0�W�>h%�����,���)�Fn�F�,��4#`�H�\�j�������U�G�j�N]q �nI�C.A��x$;Gv�]CH���7���`�j�L��(o��O8������TC�$F�br`Iw�~��#x�Qܝ���go�_h}���h�A�>�����|+?���^r��
np�>�A�[�-r�o�բa��m�����Ml���7�=K��/p}�{�d��2U�(ƴPF�1���>L��Θ�����=���0��54�W��v.D�t6�|"�E�Y�E=tA5����@y�9aNG��u����"�q��@l�)�{����	S�u1�d�2���(������)��c\�	�AE+���,�s��ץ�V����.�X_��!)l���z)a���!�������+,���{��ʟ��D	�ձ�������*���F5�]|x��jc���$�z�yar�V��=t3rH�z�n�6]�x��aU�K�ͥ���Aᳪ�U�¯��ǘ`~I�T	����n��?��Ԃc�(l;�����N���wgg�+��2�VQ�&Ŀ�V#�V�qo��W���|+�kXpE�Y1d�4���'���l�ϑ������-o'�I"��e�E�=Cq%�@f���GJbJ>��6i
B�mwx�U�������ê����X����(�!]�,%Jy�	ΣZ�鰝�O�hCo�"τ�M��H���u@��^�W���%�oSQ<9��
'�a��`��:��ЃŢ��@��a}G���Ŝw��@��� �����ٝ��ܭ�J��/����$�*��߿��_�=�JG6��^d�N��L0�̖����i:�@�gI��o���q1�d��0 0�լ����cD�-��#k�MZ���#�oI������u(0b��S����_-JJ5�p�T�% ��t��>�̢Ѝ|�%煦�h�}�=v9P��,���2����E�W�g�f��M�v���a��Y�*�E��t�Bf;2��	����},4��| d��ʑ;� �'�D��g+��+y�7o��ᦶ�{gM��W�gf�Z��[ q5hE6�X�>�Ԡ��O
	�X'���Ph8�z��k�C$���"��`���I9�ӑO�������\m�K����:A�Z�
���WU��G9a��N��"�Y����\=˯K�$? �GB�|��z��2-��P^��˗P|㴫	#��A�E�e�"�.$��2�\y�K�.ff@�ص�X�J�m�#6H� ����4�0�%��l�;�H&.�

\��T��n],/��s������Q|Zv"������G;@A�еK=��0���l`�E���S�����NTu��{V�{�@A�;�����W�7��j6�A�M�X�k��p����/�����$�IK�_4a^���`9$@є��E0nt�Av�$�3¨��6�3e�qS!ޛ}��´���ɶa���YE�
���]��ra��oAHc�ӼQ�~���;���2qh��3r�撷���<B�+�݊'03A��3A���U���e;6�Zx�"�g�my�Obĸ�
n�ru�����gMp���өQ`nl�.'���V�"jߛ�7��T�oz�c��=���c:r�Lh~����/�-~6�BNr�E#91L���>LC���M�A
֧�<V���k�U����th��\��¢��~������7H��d���,#�����b"�%*��X���?�i$�\풞��O�G�ߪ���wf�R`��r�dǽ�P�%� ���+U�Y� ���/l9��#i�4-~ق���j/bt����(�$k)�nG�5��E(�sK"ik�r�R`_�ģ�0�8�R��* ̂���N��FS�ɒ�`'�M(��TA�gt(Q��h]=�=��lUN���jv��XB��9�&z��v�Q�h�'�CzZe´��0��l�
m��ɳ%�Jah|;O5��2 ��g��<�%Qf�xe�
�ա�ֳ�X�re��!Vj��w5]u�)Ja�L?b)��:C��䃺�"���(-iV�0�ߋ/�S6�u+4n89��~�\��Ut��n�Q���5`.\R��#^��L+�.��uɾrN���)	F��f}��>\8 �8�y��r&]���b��} ��?��Ҫ5	d�(���d̒�MT� 2d!����*R@.�ۮ�5�����B���)4��<s\�6���,o��NV8i(������B�R��t�W��N�9�8�����%��T�ߵ*�rkk���n���S�nc��q���"i�s[_�<,�4;+,�����#i�u��n�R�Z�_a��8�M�m_�9xɻT�ޙӺ��Ɠ��<��d��q���dM�{���+yמ�m�7'�Σ�[lzU�]�%g�K3^�W��A�T�h[ͫ�cu��k��ۗ��ia�6��wf�4}Y�p�>5��X1�����kjr=�Y爖¤n�TA�n��P@��D���:�	���f����z�5mq m��Qz�
ͅ���61(Ha\��Mݱj�w�G�Q��y �bg�|�~��Ɲ�@�~�Tbq�]F�Z�^zk,X�T'O�r���������LL^2�g�T�$q��� M��6&C6[�t��T�9���ߚ"�m҃��{�p�ā�L���<�^Q�ـ�`�O��e�w8�Գ��X�l��NQi�@�#�H8F���ΰ��`i����hSA{�kDYG�+t�����em��I&����XNN�]�`�jK0���I�q�%�{h�T��C�Xm�Iķ@�?#y��~�s'`�?L�9���x�P")|4*3���k#�I�f��C�Пvx�����@�����j�Z��OX���Y�9����&?ȓ���e&���k�H�ߖ:��@#�.��"k�'�^�_[��\G/�k��(aag�AA^ӂ�d� ��~ގ�7�����%�݂���,dJ��-f��*����q�tpԂ���9XL���l��p�>�,_�	
F�?D�9�H�f�%�$�t}�lv��;R���-�ғP|�rH��í���I8�oO����:�����3��Q�fJ:�J �[��f%�7��J��"�O���*�,�z�������5�_�F�����37�ǒ�,eN� ��l�{T_�ØiD�Ї�*���|X?�}�ad �,�"����������_B�l|���RP2�Ŀ?e�/T����f��-�^��yh���s6�6�a�V^=�"@����&�߻- 0�Ʋ�~���U��Q+��$�
�=L�����[�5V�����,F@����9�K�C����/�9u�_?���$��8��g�=9��$`���t���j�4�)�p^T��1�j��}�1#8q��e�Nsy�����sm��'�����V/��a2KH��(��Y�֊�aſ9���x��I�����6	r�.����|���̷��p��
������œp|8���R�9�s4K�L��E%b��l���	0��@ȳ_��W������B�m݈�k�C���~[&!?-h��=1'��EHՕj=�����R��3��;0�m�%��9�G�t���T�O��G��	��H�a�TE���� ��������]��v+�$�"��x1�v���q��^���Vij��e؛}��x9�W7�IT�%�����w^S=j�=��`j�)Nf�c��Z�@%�i}z��BnNL��kpe��{:��Qk|��b�	�1b��B�=F�|A�C����s�:Eja�|m;"�]�woo����;�����M�U9�����k���>i�$�0�o
�SUn�$�U_�N���U
���ekyR
|��`J�NǤwv�fw.x�"����=+�FZKm�iG�s��oG��6��)�CԢ�\�a�dR�hT�a�ÆM��f��	'����L��W�M78��~��z<�{e3��5<WyI=0@ք0,�J�;���Aa+����&������-g�_�0)�q���Au����>���0��F/B)������2M$��n"����p�X�T���G,?H����U�\C�[�_����xm�Ţ�<�qɖ��y|U�*?k��g/]}��)�ץ�á���*��N{I���	��#���d���p�q)?7�~S��{�9��;�\�ȋ�~;�o�_�{:ɮ/L��h��&�4�t��%Q ���do��e��Ћ3=�� OA�ѓ���C�n ,�Twr�5�䣨
���v�>� ��&[��0�(n��@K�oj,�2��膝)#�|��i�ϨU�kZC�O*@�����\�o��mL7��k=s
)����P��H�&U��a����>���˳6�{?�jߞ>113�(�@��g����Z��u?��ۀ�0�b��rkS�[q�3]MC]��Ջ<��`�W�[�#��U�a�a��X��^�G�f�9ͷC�C_ݱL��;��UHg�������:F1��'�#Ra�.ܢ����9���G3����\�&��£D���zURw/�O�zKh���;֮'�ab^���x�pȴ���V�8��^^V�D	O��]s����ޖY����د�fӴ),�-�L"�o-����ݨɿ��d+�: ��P�\�VC⽼)�7*��B�8%�ª1*��	=Q�Fu{�[��´�/��;Yv)��������J��Y������{`����q�7̎s�5?ܵbz�;A\=o���h���b>_uݻ�‬��<����I(lk�$��5�=^:�����^$G�_ gg9��dl�A{U��i�5�ٜ�-�������b��L��o��0B��:]����A=,��|W�7e���W��**G�қ9M�zsZG7�5�m �&O�e���,+j�ݯEi��`%Bg��N�������9:�>ٶ���6rt����=�7�ᕮk�=������`�ْ�����Ϭxm����a�\�\�h�IË��_iÃ�A��%�Q�>2����o�'��:V�ytx�Z��!D�3f�(A��Q�U�1R��cH�َ�t(*�1��~]ȹk��ֿ$�B��Nk[��-O�Cl���b>������C�m�`�0��L��7dl_�ȱ�I�	���%�Wώq��4�,�A/g�!��zι\�B�6�6\g1�)#�a���������Ec��}_b���*�6�L�i��B]��ii�J̀&rn���+�@�k�GkGՙ����7�g�5j:����� �5�L����(gL@9����9�<�DQ�3�0i'^)"r�c����� :c�{�ܻi��bm����si����Q�f�AF�����KH�d�ϭ��si���$y�Q0����#��'���%�#�@�c�TM������/��vQPe)qZ��#���ƽL�|N_eiGq�i]����n=�QZ��,��<5�}I�t䑖���;i��ٷ�/���əp,�2���xXlxVHYEB    a482     f40U�;GvvF�P`�i<�$ڛ�,�jt����G��*�͛�7x��0eM"��V�����XB4½?�"���!��}Ȕ����������K���Y�����:��M7�Dc�����z�7�<�+`'�u�X���_��?������߻�KϢ�k���XÅd�s(�L0��K��$����q!AɩZ��!Ǝ�Z�O ��.?���h�a1�ȯ�9綠���"޳G��<Y��<��ı��JB!�8{Z��i�跨�[�l��'�Nf8Ҥ&%�߲�->j�.���U���Nݣ�[Zs]S�1KT�d⅓fk*�u�lu{p�B2<M����g��(�W�1������Wf�0u9Dk��8X���ә��ON4ɱ�)hw>�l`�%D��.E��P�Z�����m�@VS�/b�ȣf�(�R��C��[�P
�[a�r�/ѓGS�5�5�1L���cm�)W�{�=n�)���Q��n�q'c����^�$��J_��w�R=��l�e�����/{���O�"���� ��t9�������򼈞Q�ܬR�w?��q�e/�9�>���a˝ł͟���>�B�8�UK�����-���f1��I�)�	W�B;�.��%�Fw]��d�O�V*���4(i=�i�G���)-Jx#J��
�+y\n0���d��.��	-�6�C�*15�_*�Hw!߫�y<���o-#I䣢d���J���\�Ru��2m`�w� 5U����,AGj��l����0jSF��mW|��[��PqߠL)ϝA�B�X��k����њ�}+�����JΔ=x�=�zME��w��6�l-�[{(��A��pOX�즱�#^�j5j���Eq)R���z@?�T �w J��W�?p�� |T��L��9p:`�3E~k�\E�2�����=Vdvz	�̄�/R�4⋠�B�%rac�aی_��J&�jb�ǊJef9m�#���ɰ8���)���/�IV�f|�q8�
�,��p�n�����e)e��EǷ��r�;�,-������:��� �>���=(:z�����@F���W1�xS,3�	G+j��?r�q��������g�!\2��1^����͛6E+�~z*��=�?6�tZ�O��O��XBM�~7�Ep`	kYhi�����s�K�sn!#N�m�93S%'<4޹5���4�_m�(S���U���-��ȫ�=į�KV2���H�@�"q�Y���-R��ė�p�����?��7��]W$:.��;e
�G^?�m�Y~�g�+��G�
O��s��\!��j#Y��kv�ĳ� ��,%_bwp�j��%��hX�9�O�ًx�ib�q.���=ɀf���j��}.�6�_��m4˞:�e��s�ɷ��]�.9��rq1!�]��b�z��ןX�H/v��Y�������X!jn׵Q�P��M�T���d	ւ?���no/�h�	sI�e�:��fm�?�8v�#6_�x��Ӣ�E��n�m_r��<�i��AW�MP����m�Ix��>ݭv���$�����`��kh12B���x�3�"�O��~��j��a���kE\D;�ĩ~��q,
��3���F�|K�����ӛbi�y�� ��AW1�˃�Au!.������B��7�6�����Y
�Id��M�)ۥr=����b�xQ>��$����\��&� ߶�T�^wԕNg&�舰F�q�����!ڧ{Yq�`=fG̭�WU�K��4���q��V��8�~ݝ���n�}�.㝻�A����9O.|e��-!���e�W^o��3r�����-`X8ر�N]�-͒ �UA����Nl!Mx��g���X����n���X�K����c��@2�����yv#�o���7V�sп>�d��I�Iû����OQ���<^�c`����V|��t�w)g�����=%!}��F�tX��Zc�W�ܫ`���k^���a�*��fej�+Q�����;,!І�}Y;'VY~#5����8�O��Ȣ�����Xnm
N�Ş:f!���7���i%�}Ee�˅�1�GhȤ�.)��'�j������ *���$	�������0��]J�i:�@�5�(�9J!��;�yb��P��E���t&\3 �p#_���I�g������c/g�]y����W����rj�����/�ck.ȔV��}R�)��$�^�@��1�|�� A�ʯDB�<�Y�>F�t*�O�JK'd�����<�
'���{2�z�����j=�Jcpu�7�i�/�v�ΒW�jJ�n����F�Uӊ��;��Wv)@��Y��]���w@1Iw���"�ݺ��č�)uHy�e��Z �1t��s����	�5gU��[���^�]�Ӌ���S��LuE�`-�Ό����W����B�v�3�<ׄ�N�# �Z|�e�z&;�+�����_Oy�����8B~�be��Y6��-�ǋ��A��X�zf�����Ev+R���U���	 O��??f|y ��8���xIZФ��k�����h��͒���|�����L��I�%~�k}�(�$�B!��赂�<nҹSU�������:@?c�-{�M�2AAՒ���� N�9�N
����8o�N>�������A�L����1��f�_��hͷВ@�f+_�D!��� n�5�4�2�	�x��N��Q�C����q��m�����,'X�����r�� �.)�V�^i���q��`���;t�b�_�8�'�KJ��w��#uGHh���Pf��x�eesZ�X��y"D�`(R����k��t!�i�\�=�4���%����mqR�L�[.%�4��%�g��Z�N��s�M$t:�&�mF����K��E[wl��0�;+�L�W)<ټ�w�>ĺ�{oKپϬ�O�{;�^���z�υ������U� �_�'Xb{| [cv��*��$���W���^pW��W�{K�B����T�z!2y}N��do��~��͍%K�"օ�� ��NP���TRޅλO[t�Of{���A�"W
�|82�V�gO�r�4�Z�o��$Yy)~'�ҹ,���;��x80�:�o�T �����f�I��KR�����'.2O1,��؎��WEwU��<���>do�Hj�AVA|߮���hYѢ�s��8�����C��)l��4��^>1����op*L��i/�*�Ő����r�֍��?='�L�Z_;��oٵ9`šUjx�ƃ�n�b\��0B��:vѩ��^;�D�k�7�Ӣ̛���A}�i�L��v#��֐���J&M!:��ƝBy�3���~^9���݉-��6_�͡@FV�:�S��/�����}ֲ�of)ʧ)�S��k���M��"pؽ��Ǭ�O�S���3vJ���������kr	xw(�ѥ~h4pT�u0K�D�^s^�Fܠ�X��ƒ4����u�F�j��7)��~��)`�cR����|����(��\�Sۋd`^�*����R��6�
���.��K����1q�������0�~���O��W���y�����H�zƸ)�[ I���J"#�~b���1hd��������-IQ��j
���}���<���B�7�6��A�s3�\&�������ߊ�ꭏ�^��'�-��[К\���(B*��~�n��iB��/�T����%�(�9�e0X4TOtpj6j�U�_����&ZʙJ�`���?|B�"�*���x�✿��K�$o��_v�(����xerD%���:^�߬0�&�eڢ�p[2�n�����"�]��f��R�l;�Y�MP@���;]%