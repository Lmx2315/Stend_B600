XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����U'ڹA�I ��S>{��=�����&z4�7�<�z�lL<\��B8�(%
�����Rg@���7�����\�����ߟ�����gT�����Vw�W�����)3�V�Hm�:�j�p�k��"�����K H��x%k�v}Z��C3Vc9>';���[���C��=�qayF��m@֯L��5�)�Կy�@�q�	������޿Y�ޭ@3$'�6~�@���b�k���~�4#޻�
�u�ω�����(���3vi)[�u��=\%>��%�mu$G�6�F.�:ӷ 4x>`L��J�� ����X�T�&���T����~=��.U�{��o���z�;��b/�ˢ
��+S�tGO*����8nL�?�g��=����v��[{��S_��Ŋ�%�� M��o��3P�������Y�>ՏS��?=�����j�r1|g�C�-�\Ψ}m���}a,�K�>[����k���c�Þ��6	wև�qz��޲O9C-�E��J	�6T[�#�ڌ����r��Ǯe#�Yhӏ�Ǘ���~�!y�&���;�WI�i�u�&���A��mt�~0bIL��6.����4[���F�/�<��
�CSg����P
/d��Ʉ`P�*�uͰՑ�x'�e�.Tu���	���n�l�0���d�D-��P�����`�o5!���ٝ����2�E �L~{p{����_�'B	�����A(k����D��3Cx�&#�:�IXlxVHYEB    11e4     520'#��yW���{�))ν�����0���7/p��l�ۺJ ��V�Զ�څ����tH�.uN��L�Q���m�(w�N�}�!�������r��
���w4��g��^O��ѧ�v�)������{YI���D;�8TB�T�]��J��[k��1,��7�M�P�|*U�NH
{Ϙ�:?���\:2���dNJ�%��1�����7t�(�W3DУ����PN�;��m��Arc�eJ��ĔYb���`G���Xx��]��VT��Ӎ���$����b�Fs-�������-�|�$P�*�LT2ȭ
��,!��݄W����a��ERK��F��45�ȗ��8��n��&K��Q��ᖬ��%������1�"ZO�;�����OL ']q)��9�`�O+q��)�[�t��V�ݾ{�n��&�7��(/	�������8�{4��l3D�º�#�ru�N�g�_@)�4�!�KK������VP��� ����F�}ע|����V	ul�kX�I�9w�"���[��Ḋ��$b?�]3���,�M���gx!�M�6�@ok��>��)�V�%�`�f�/>��Q�aʗe<"��]�0�W�d�DJ�QI�2�"!��[&�$-���Ϙ�L�Iw�,���p)M�־<خ�G��oML?��;,踊�V����$/B2��on%���H"�."bp�|H��-���v$��q��9�/�\�0��xk��nr�J��A���%:-�ճ%���$o<�m��O�1~�N�"�Q�x҂�bH>���	ƀ����D���e��!�޽ID,�A�z�<~�`?�
��J ���3U�|��!5}��mo�O�8T��/�.�T�|����?�dx �
v����֠�E��-N[1{���z���`�%�_A)}g���)�B;(�� *�m��"��5���N�~��tm�G�ei��I�ވ��ys`��{v�Dm4��J��4�M��<�����f��줒J��V;w������9�h�uO�M��������~e���u�z'>f�M�n��p�| �7Qq�{s%�F�,��t�#v�_Q���۴_nc}�l��{Y��x�
w[/�>J?�Q`a�jyH9'��Q�ϯ1�� [��cr_��P� a�"4(4���N��,�m�6&do�;���X5�&��Bm/K�G�u#���20�+J� �%�k"�q��D}jNV�zU~O�^�P��%��G];�6�a)��Y<�*:T�Qe�#�f�G(��U9�R
~�(�a�k����