XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����6���>M�37N���~�m��e
��c��PG;�Tj�s�a�_i9�\oT.����.�.������ܮ4��Ϳ]��{�Y(�n���:CP����=��2�d�l��}&Q
�[��č
�_�a����K�D-�84y���������nq���t�9���=r��P[$�U�Oig�"g�u6fY�>��}����������k�h�\�f������ҕ�޽����@�A��4�E��.ʬ��4Y�.�Af(��c�8D�4O�oMvx���η�Q�|㕲�~v�,�N �g� V �� V���"oy4��py���jvʊe6ت����24�=0�+s�;�v`~xT�����6�*<�\�����l�h��K����><��&A2��=7���L�&�ZT�}�j"��Wº$��6�f����.�K�Ve3�b�T�G�V�%|����9�oߓ��**Kش8ho�.2����D�
���͓M��ʞIh��gC�փ���k�Yƨ4�o��H'B�+P�xo�񽣅}QCOx+'��=�@(QŃ����t�W�h���7��̹ԡN`d�,Q�S\KP������ql��=vh=Kv�t�M�T�)��ާ�� ~ĸ�� �k;�jـ��<׬�r�v�>㷄nZ�fؚ��aMh�Ꚗߒ�$J��]�F�9�C6�nK+|�G!9���.4 �A�h?�"q��]c�t�D��u�>[+j<f\�g�;��9��7���w�XlxVHYEB     7b8     2a0�c�I
�s#3�T�#X����v0fEh��3d�"o���5-��^/�םh651!M�;Vw���_��g G�)�9��ŔS��&�B�Tp�>a5�11�ϓ����=>M#��4
ހ�ô�:+�LK%Y�X5�r=vσy�2���t��	�+���T��bJ��jf t�Qь���A��l����)�rY�H�x��2s����v1�/�3X�"�F�'��<�]��؝��(���=���u.��kY*�%o#�?ѱ1`���� �$�'+�gq,v�m�Դ���"�� +.\��;�%��9uН]�+�r@V���Hm��e
��!{j��
��j�M��	
����J��CĊ�R�����wU���.�I6�#�*���4_=cŇj�#�W�}�ew�B!o���%�X2Pӕa�z���⍯�i�m��ɇ^ϯ���NdZ>V�8�f،�N��$�F��Z"�:�x�Va�m_B�Nb�s�#��A�co���<	D1�FA>�bj�ȧ�ZnÞ�]�r,A�2�Y�,�X0�����on/�A���vz��y[C��=�=eS�����]����ќ�,j�^�X:p�Xi��ΜV���I|mm����8��~ݱoщ�?��Q�C���b�,"��?�4>�W�3k	J�3[;�˖����v]*Vf