XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������x5�'���Q_<��m"R�]�\dlE�W����S���7�䥈)�?	���`�GUކ�^J�a�ﺷ�d� ���)��L�TE����#�����F��g"����N��DK�	�=�U����DN=������S.��� ��T��m|h����~^D��j>�Q%M���@j���cm�h�X*�c���!Y��)P�}_�QV<T
X ��oQ�p!/�	֑��9E�0cS[x�v/�||�4�������Z=XU�&��\��sjيaF�O���]IwoԿ�S���EЊ�!�;��T�BKC��*3���R��4�$Tk�M;�;��vϕN'%w����4ķ4M�cY]͢Rf��1�Ru)�	b��럇�aaR�+z@zS
���Du��G�I���s��pi�^��h�H���0���K�M��,0�j2�L�>q~�r�d쐌���{�>����H��م9��� �`��4���vw=Umk��� K���Z�K����"�a��Z��8��s����F1�F[���}���O�	�AY�@X�:.ܢ��j��&x��2�͐�2����~o�C��s�,5���uFH�J��庪C�c��[�r�+���da��I{�C?���5	cApl����-$�a���G҅H-�,�C�\(H�������x��ƺ�� +����,���p��wy� xO�xS������U�\?5.0�ţ
�N�u�]k�T�S�#����XlxVHYEB    1047     4a0VXV���	�嘜=lͩ��W���e%���N�Y���<
Q�A��ξDC�Z\�s�Z B��+?�M�F �尳e�7�:�2�Z;���&����#[8�I�U�S��l�jI���2vy�[�+n.A��
�L�)u�Xdm�th�Y��-��T��s��K��V���Ѯ�M���Ý u�.��6�.L�����9E�Q�L�"5 I-E}�*%:`���6����I;4C*]�T��H������
�`�jf���
�Ϲ����bͶ��#:��QLQ��8���P���AC���uj���T|V�6�C�o��^�� ��|kV"P�
�[�\:�i6�s!�YfC	���4��Y�d�u��X6-��gl�m1r�kkF�_P=��6�+�����_�g)� �a��e=�ᨔ�{���I/�&9K@;PA�9ϕ�x�%vJ�^�8��^/>������5�@�_�q��ꐪYwd��	���>_A��XpI��O�1D2�z(;�T)ފ&0��[�T�C��^|	i�U��t?= E�u��\��MHx-�]����7�v�W��0������ٱB�O��#���G��ӊ=1�ԍok����F��t����ca
�V:�ja}G����zg�`lݾȻ�2�/	aU«�'b-����Nr�R� {uW��x���?����v��X��)@ �V���o�'�h�VB9CQ�X�dJU�J�*RK94�i���T	"�x�����dX��ey�E���A�=��X� ��k����2��NB����8RCR�B��*㖆Gճ�d�C�AYۧ ���5��z�&f��bbZ
���\5H��9�(�������!���:��}"s܀`zz�W�����G�ȸ�=����p�)��"+ ����4��b)��)8�����-�\���|���e���a�������' .M�����l=�b&� 텒i��3T�	bS_Zox����D��2�.�f�h$��Tx���""�L���Y�w3J�C��q����`��!������t���灃h�'�zH�D��֧>�#������4,�:OƐaQ�>��C��Dm-p�>��ު���	 �;�p-�^A�g�h��i`��n�Ⰿ��L�f�-�S����)�����͘���R\�ܖ