XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���"H\}^92��
��qO��1����ГBZ
_���f)�oLpډ�)�5>Κ��1(��T�"��,�}�T�U�a_���^�/*  .o��`F ���e 5�|��D�Ә�$�)a_�ό���o����"��0r�m
�$��a�#�ТG�?��0��gJ�+v��C������"#X�Ҡ�=�8���Ķ{xp#��;��Cv�7�`D]�����e�uUw�a�I^�|9f`�3�n0�/�F�Bh�u�U��(����WԶ���&	)nϬY�-0�#&������1i���u��q?�<�YԷ�\���o�R~PC��)�%�fSG��;���=)��M�L���@��
��L�������-�a1h�=��T[,H)����2�Ѫ�v�fESG�0��Օ�?��O��	ҔB�⭸,r&̸�5���I�j"t����<��l��F4��O�`-��4U;i��/�j��0(���Ժy�7��j��r����s�e���S{�zۤ�T�k�
��sS%B���*��z��ٍrU��&j<�?_�����e<��Ao��u��M}I\ds��T���Ac@�/|_� A���Ԁ�	�ՐA����!S�N�T�
�Pw�\��Ņ4���,g������TZg�҇5��i�T&Ԍ�.O_�f��-����!���|���4�/HWѧ��$�K����CE���;�U�v�ڕ�����o6?mjUW�/	���&�ޠ��U�{qݹ��XlxVHYEB    152b     580b3Έ�='�h��)G�I�#�a��4�����B~"{��5�v����R�^`���=#�;��%t��p̄)�j+6�����3Y�5��vȪV��
R�c瀜%�Ӫr#'Y7��$���%ϣ	C�嶡�Dȶ�1��C6�<C��'�"pɿCr�]
W���c���.�DQw��$�q�ۮic��x��=�i#\J��D-;]U>�؋sw����ؒ�I���xU��"lu�E�:z��� ���V����h�R�pwV�0xr��a��~�����*�O�d#�KN+xw��e���U�T�R��[5]�E>���|����޻k-�J���S���i�AGi�2�Ñ{+�QEU�nm���0f�F'~�KD�	�T-��������{';����;��G��&Q�q��+����QX��c� u-H��E){M�LR�;N�
SEϺ� ��l�"���>�p[Hi�E/�}mrE�g��}8<�c�uiY�-�E3�D#qh�n&���si9�a�?_�\��fT�}!�o��|�g�.ןO���`�s�Zm��2
�♱�k�OABZ�Y�~|k�F�<�;�P��ֳO���G &��4&rBz���Oj�M)��u��B&���iI�ɧ�y>�x�)Edx���!�Y��$ޥ�ET���j.I8��Hi��{iq��B�����w��"^v0P7r����9+�U�v�y�X6B��*���|�)�z��pI#��E�g
V��+�ƥߛN��:��Bs�׽�	 5$��H���l1={Y��pW���!9���o�-IG�	=?�ށ"b���n~��ps����2�����z��=sK+��ԽWxK.#IBtE4}�~����yؽ�e�']�4ˍi~2��<�nFb��}4a+߀RTj=Zz��,�i���ya���̛t'XkD���"5`LNo�M�]Q>uٓ����R��*��=���h@����>G�z��/M��sҾ���/�QȌ
�s�`�v���?"[Ǿ�T�h8��:�P"�2	\^y��zk�˭~�{��>p������Ad DC�e\7���pc�N�˹AX��}����n;Uc�[L/��[��=Aj���N��Z,3�6�RB,�J��2j|nn#_�J�Yy�_YDj�� %>��+P����v�B�-�7�ZEM��� p��Lxq��~]_c�5"k�ŠBD��v=.���vhŵ�s�!��j&������U�ٱ���1
�c��4m
��C��������Z@ ��t<�(�wX��X�O�D�B��H�}_���?NU����x�ѝm=��ݜ:&
��IE��*\�˂]P�
�0`XU����_c�j��bf`S^/��U��>&k��pC5a8�V��$GX(�K	
��Y�