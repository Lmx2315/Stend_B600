XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���t�9#;$j�В!	V�9gm�l���z�@!;9h'iS��VϞ�l,1ͭ�h0~�����������yaT?9�y������?7��$(�H���ep�x�;�����B3&L��wc-���畢����Aq(!256�a��v��׋K_*�ݐt��{��.r]:� �d�t��O�Ը��� ��p�x<3́c���u��
�/��-��81w�I-ܺә��П����}��ksk7��+��̮#���Ff,��D��A߭����/���lV2L�k��l���m�>��Q#�!�ًSqM�_%�Mv�ꥁ�F�p�ݸ��e�x��Ћ� ������S����������\�	�dݡ���c@%�jA�*X�+<��W�j��d�Xv�΄����V����bΑ�+���F���o����C�8ц�WdFS<�Os�A����Jp��!�n�Ti���X&ҟCbi�:_+ad_�fz��Ct�[U�xM-,�vn�������T9�e�hs5�ʆ��=��-���*��v����޴2o����#�R*߆�4�`b���jdS���M�����3	���s����Nf�Q��HL�������D�A��Ί5�z��~���v!NA���E|
�1HS�9��>��=���|�_��H5�}�YpM�&�K�k���w���KIL�X�i�݆�Vf0 x�ة�yЙ���������yu;���`,Z��|S�]�2�+����-L��Q������XlxVHYEB    38f0     d30�>��r�2�Ԗj�bY���5a��D��!�m,eI_VÜ��ܖw�b���YS����d��dr�>�2��<�oG����q�t�������ZS|� �D�_O�����s�f��e��|�|�6�6�쑁�N���O\&<

p�_�k�J{�rvw
�}'�ɕ�h^�IjX���F8PG�"�PK��J��藠a|���Ws灚[���=��v�g��P�����	="Dsw�H#��3{GU���
�C$��A��A�!3��j�2'r���歒���@�4���vW��RCէ�&3A��%�X; �h}�-�,sbt�xx��7V�޼�ތ�͇Y��n">-uVZ���o����۟r�0Tk�\c�/��H�[�n5�^�[f8�����8�몲�~te�x�kv�o2k�q��u�n�Ѳ+k��ٰ �"b$���m�x0��4�d�+��쫚d��m!Ե�Ä����m�^ܰ׸S�wo����q�cO�0a��{�vg�ɜ���唼�� ���?�/��!G�@�:�$��m�22���� :��|��6�'�����%��Ӄ��>TOo���S��z2�~�i@4����LͶd*�����|ۭ@�*�X!��QOu=�E���x���0�㔤֊�R��J�?	-v��(�l�ӳ��vF�!ڠ���(��H+�'�<�/�n���@h�9���hx��ʙ߷hÌ9N��9r�h���f$�������Ũ3�� x���`w��37o*� 0����JL�KL�{/����n��$u�(��QLۭQmC2HK �t��EtR��[=�l�dC�zy@d���*fņ���/Y�[9����ɤ��,4f���X�6P��zs�:{+�-�ͫ7�ݩ�:���3�&F���GTy��I A�ek��X�PW�^����ͺЛz�A�ZW�ج}8i��&��D��7�
����/��5)l��<+f�B	��"s�YuT��mjE�S���{����6�zZ�� d�HK�g]۴�.��%���[����T�v�>ly��f4M�EROV�lwY�.�����rP��}<�Z(�y#���Fp��y���xR<n�� �ʅz�V���lM�����3�I	k:�n>�4��c�ޗ8��"���}���{�y�[N9�C�N����X�7g�4m��"��h�i������x�rh����ah��_�	=>������_�;��#]���u�a�z�����U�$��2՞.�^V�u(���O����s4�ʱ3s�*;<��}�N���,lw��܇L5]�M"3�]��	L�ϡ���Glo.~��fb3qv�CL;G�Nhھ��`�v���7;}�Jd�������8�s(6]�ʮ1��7us�@&wKs��r�Ӽ�0{֓p��O)�.�{p�*�C`���;�d�[ah�n׉����4=�51�/f�	�*YC�.ɚ��I��w���\F�}�Ī�IB�� �jU>c @[���������#s:�ޥ�Lv��l���E h}N���gh�L���\��8ǿ� +	V�yK����?�������D5�������f���U-+��c�T2��H��A2�TD��C������!�s`����Rؕ-1N�4�P6�ƃh��UKd5��|� 7��m�g9��6���5���~e����l�ݗک�qCiuyd�L�h7���0s�Qp]cx�ФW3Ϗ��E�#�(nΪ���~��C-Z�Ѹ��Քt�v�!�v5�:��ea
�ra�CpScO�,uY8?# Q�Y�����#��~�0A� �M _�/"V��A����uK�|mg��7g����|��{1����	������Z�r
y��2fދ3k�A���z�֧�d�0^g\��pSyY~�e|��Z/&�%5ʷH����,h^�y����L88!�Cs*`�_Bɏo��3�`T2��rtq~�+z'õ����E���<��%�	I��2�ґ�ȑ�~R��;Y��Uj�%�i�L_���6�C��q�Kh8P�6\]1߮�څ_�-�AGH��*$��ҙU����T~��L�>��I�TR�޴�WO���w�8�%ݴF�Q��gh�qx`!��m=�rQi�C"(
4��W�� ,h�v~�um�_!�#ղC�q��ٍ2Ǽ�Q�7��ն�8y+��IoH��|QyBNL���Y�?�]5Z��p	?ŝ���2�lq���>.�Ɛ7 x.�OA����>�DX�g��͝��o~����]5���ݏ�n�	�VE=OT�z�v���r�҉��"+�_>��A!el��ؾ��98E>�1s����L�Ȣ9�c�p��H�517C����U�~))n�Z���e�ُ�ö�j�C&�����$�g �-���B_�[����Oz�ac
xaUE=2�����Э$!��p�ς��8~J�|q�ل�["Ơ^��c�#L�iő�e�o9K�E�|f��V��E���m���:kf��춦�A�Lm�6?� ���|���hծ�&���C�2�����~�]���5�o�� ����P�@`WM��^'��}�C���)!@"ٲa*�1��9�T���s�KIۉ٘CӺ������������a�y��hJя�;}��)���҂ˇ�<��"��A����'R�6�h��w���{��JSP.�0�ٖ�'���W ����8̯:7�ER���S�8'n�a�(��� Z���>�gK�Tn49�u��bku4M->5���1��TMG�[��S�e�Ċ��a�2����+0�4ʙEǴ��S#��[#Ó�>��g{^)ψ�4Cڔ6j�Pt$^�jm&� �� ������ފ-�/ L����@��q_�~e��Y!�o9�[�0떠P���&�ԋ�'r��v*Ձ����zD�	!�_��=�������Y �FN��Q��N���U�>ė������v���w<�Y1���~F/F�Atؐ������Yt�`��kBy8žFP%�;��d=
�N��B~�Li�Xzx�r�N'Z�l
��+�E6:ǖ�_kUDGuI6֖K40'Wh��e�,v�vIH�N�rC�m�l4�,��B�w(�Er�z��g(� 3�&j]���H_�_~v�K����������h�G�'��<��R��e�es  ��q�A�(�|h�n�w�̑-j���RO���`]�i/�����:��mBԿ�ң��g��8M,̟,�>����I��|=�<^6� �|ʆ��1�n�/�+Z��m�%yNiX�RY�T�����sy���4��|��=���w��&������4��X�2��%-,Rُ