XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��/�8x*��P�J1���A4�(�g�Ƿ�0�����w�ov$=»�k�#�0�.{$[ų��)^d���+�Է�EB�t�c9=H1���e������T)��q�>K�jb�~#�\P�8����)�S��7A� =$i+�ww�J<�~��膯p��Q�JDr��T�@����Z�O�j��%*\��ՓǿKY��0��=ƹ=^��yZߙ�H��j��^�
�˯���RB�%�Ԅ�~}\f���ڔ��YеEif��ݧYh	ѻ��"6�TA�vXU�d}&��.�`������1V�#����|�
k>�0#�I& 1��?�G�gF�����3N�:18	e1�%>� !@ύ�Z/	:Ğ��n�7�.3+*��=�eq[T6e�$0�_���b����nx��nZ8�ʚ��I=3�zd�}>�zV{1�v^~�P�����M���v�/\�OCQ�S��)�c�#%K^���:��!��q�7��ǿ3h Y�Mc�K
��œdQ�yX:���zB�%�8gAc�>�gK�c}�,*�0�XU_K?���	�ۣ���A�'��]�J�d���������U��f]�q3<�IKB���j
��?��J��^�W�Z??+�c8��! w�;%68�������>E�O^�*����8�������6�J��]�nB�g�)�~d�*�Ѓ�+1��r��P�2������A"[-J�ߖk ���R�~4�W� �5f��jC�["�����l��@R�T�s���Y�ɀ�XlxVHYEB    7945     7a0E]V��%��jHA�$��@�X3\��e�J�v��w��JZ-�AUX0	t�����H���#O�)��y��d���[�Bb�@&�U�<��m/X��D�('�Џ���-&�v�橨rc��N�ވ�%jZ��du��O�X�w'z�4qئ!�E�:�¤Z��Jݼ00����Z��"�c/�|i1�׳����^[��0��Q/�Lˎ����O1�O�6��˜�Kأ^�fv3��I��C���et�oș�:�e����Y&!��C���f2���[]�=�ߢ�=Dν����F �[�{&�W��%-A��ɸI豁���TM-J���{��n4ph4��Wy~��;��{ڇ'Z���)m:��٭~����س����kVߺ��hZ�/)G5�a7ys�|��xI��x� ��9~(�T�y�Vt����B�������O�>�E_.P]n*F������=}�q�G 9Eå�K�(�������w���"�{Z �����ʜ�N%VQEހWV'M�sf�#�:;�����#��;�ݴ��:�@-��8��!�`�t+��Q�S��'y�n����3�;�	�c3��)�������%����FXN��`0%GuA����V���P�)�(��ϩpr �U�C^��i�����OA;,Ӗp�F�@�W�´�4��YXC)?�G�j<�Y�W��a?�AA>����a�!�"�˾V�J�&�;���&f(#��G��ӎ���S$d/��ɨ�+�.`)]pa��hyd�yvk�l����{��UJ���8��s��0�R�U��3�#�N:�n»&���Zl��N	P[� +��8(R�P"�ίw,���w�0*SqP��K;@��Y����s^��؃���D?�.�/��X�7�����7���r�L��e���`snuwp>�,��wi _�D�WP���Ф�x�D�����lK"p��i[�6���E�=����S�%(��V=�O�Y�/��Xy����2ޚ�=t�%�?H%m/��.Z�,~�F�Qx5G����n��/Wk�~[�:{��௤"�y*`nh� ������o�E/Ra�9�WK8�`���(�q �D��x!Z5Vm=`q/x@�h-�w_�j/����VJ��YV���5��0�B53�9:��*�]N����r-���~BJ\�D 0�|����m9�a�75V�^%�G|!�7F�*�h<�ޣ�3>�\g�n/��J����U�8`���`|�
Z7y��/Vށ��Q��]��&+E�@��j�Aud�s43`4�t�����
	R����[`�{\ߙaE�Ե���*������Zw�'�U+�b�"Oޜ�:q�o��[����َ�`�o��������'�D�F��z9����":��
n��HC�k]�'�<uV�T�^9TaR��)\�+Ƚ�[n��.�ϯ:�r��?]݉��ٞf��	���
.p1�5�A	ꑗ)m�eA�JU���eJs�7�Q�<�T�M�3��擄��f���,aYRH׮*Y�E��8�W�����Rr��Sc���쫆c��%0qͤ����F4k��LWb��r�B�hJ�ƚ}��xU��%;��ʊm,1E��#	x��U��#P{!�OT�C�{��f�����'�XI�� ��P���4yAD+��Ql���TN�c�8+`�7�M�ķ�e�hJ�������dd�<�Sq�3+����s���7�k�rn�z��2����ΰ⨥���4�t4�3��ß���<����[��}wv��I~�g��fR\_y�Ƥ��N�t�,rn�{�������8�o)u���ϣ�P2#���?iNI0�У�ɚCl��LX�H �����q� ���ĥ��wD�P͓�1��z>����v�($ͮ[������ߨ!`�Y�9� y