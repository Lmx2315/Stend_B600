XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����5!�D�$yb{ād �C�zZ��y�ᇹ��D�pQ𗗩�*�,C��簋�Tn���>|yV�����5��h�'R��2Q�-�lk#�~^���1�U�Ft7U�|Ƨ�ހ�V�6�!��̵d+�,�P�2I�?7�ej'(��@3��|���>�l�r!9��/&�cΑ��T��_wZ�{	�8ȝ�t	�j[�jj�ѝHO�}��
���@32܆���=�-��PfT�rO�Us�9P�8�TL��>5��ۺ�����h��ֱYe��w���}�]�徭-j۱�Cنb��;í���Q�i|?�\�)��~.y�ޣ�Y�#��*�K(��>$�@�r�Ⱡ��D7Q��6�@_��n����T
co�
A-r�1��r"��	�<�?DY|B$�?�BC���܎�k������wiZ�钻M�e�[�%�ǻ�d���l-�P�z9H���r�]��rg  E񐎢*�(����nqN�d��?�y̏���}Ÿ�>+Iϰl��:"�{��V�G���9�U�(���}'S���9Ub����T�C �����7ߠ�!Ƨ��؛��KHH�����ތlV�v�ɰw��fS<��`�	u�	��Z H��(cɁ������Lb�:�t�c��B������V�:oRk���q�GD��稔�榚����� �[�D��h���H��~
�!����4A�4��%�gq� ���+���Ւ��p�d<�b�0c����}/��TJ���Y�ػZ�h����F�!xXlxVHYEB    8625     ee0K�4�<}:7I��M�u����rJU71�n�S�L��y|upj���O]�s���w�G�`�D~j�Ǖ�w�?�����,�`oE����4���P��kV��%5�(�#�����Q�U F�r'�Đ�;������T����r�Q/%&"��j�ƒS�������}x-%���P)�	�B�������Kׅ�b�#�f�Ԙª��O�s����F���ޓ��a��p2�G�!^�:3��K�F1q��!��_���k���{qub}���1��5h�q���n�Rx�m�� 4��r��&�F�A�6R�٩f�"��c˲Oõ�c���/�zl��&R!L�*�B:��D�'����$EA2��<�']1H:���Ӊz(���8�u
"��b ڞ���nP�k[�7�Ș��h�EN�En:Z� #�s!%��ˌw}Wa�2"�3(A"�A˧}��N�T���V�$.�4�$��������x����د��|U��0��X�{˭-MPH�Þ=1D(�
ԋ�;�4�E{��?gy��9��V�p ���H`m�$��dF����#O�{f��w�ᘻ�3��Ys#��%�Na};j��a���^�0+� a�=�#��:��(+s+n���8�Ղ��R�t�V�E�K�6�M��E�W�;��+M�A�(���Nƨ�o󌲁�����6�S���iPZ��{���3Hf��M�k�먪
z�DT��K�;�
�!9�6��K��	�lǨ�[��)߹]�=&Բ�P���%+/g�1�Rr���!����ĳ��CB�:��K��ou�_��e����8�Aa�
)�Iv]3�ݒ���$��T�a*���(��=�>D�@k��cx�b�M�2�3Tn/o��x�����B���	Ќ���`���As��ўԱ�Xt��n7|�I���z�؍u�ɘ������>�n+��ZJ��Jx��g�8dk�
�$�x2�	u�=�s3�(���|#����<�(�&u�H��Kp�<��P�����DU����>${���ܑx�O��[v@���s�q�q���k��]��l�u�=�y�\SL���}I��&W��+͹����%ً�t��u
��%�%���KN�"�_�;2I�{sx[8�g�sJ��rj�E�frКҴ��@���`'��կ�c�M�U���FiSx���	n[��B�X��w�dr�7������tU����l��P�;J��X$�_�plx��b:�"�U�"��8�ݪ$������wn�fV��nŅj�tR�E�wS�6%lO��Ă:4r�JF�.�D��U�����̍mB�:�5G�ȑI�T/�}t
r����pƨ���+ъ�1���X{�m�Q�[�Q�KO5��������J�uSafq��YC.]���ޮ;��b�,YM��i����|B2���ʛ]^)���[��P�ez����C145 �LhV#͚����~J u� �1x�Ɲ7�c��X�-�3�I]-?�-��h���ܑl�_��D�$P�2�Ӫ0�W�Vw#�6�d�02���N���	uERh����
��=���gsv;�ьY��Q)m�|��e���}MğL��G&?���xU�p�Ӎ�S�VPg}waZ`��a���I;$ ��N���	�r��M<��3&?�]f�'3�{hs:Z1���N���۠&���9ǤԻ�L'Wh�i�0����Y�)��c�%����Zp2;�����ݏÉ���E b͆�!�=T*�ީ��A��:�[N��m~|�XtL�{A���6B�h"��S�|��n4fm���P{t*��h��Ln���kKR��K�E���DVU$2F��N�OxE����xF7����TjAO��[��o�"L���*ly�� ��d���� 'v�b�VOq�u9�ȟg��Z/�E.��oR���0icZ��� ��Ї5ۨ�%zT�Ѹ�n�$�QG��Y\�u�'zKYX%\�#�N7�_R�;�*R� �rօr��&�ڑM����"")k��}�ABa�݋
������[�PH�O�1/%3��v����P�_ʘ B.l�
&K狅�P�4|�ϡφ�c9Uܒl~Qm��(����O��c�g
���w�#༗�j6U���V�.�2�S��]f�9�J1p�rTT���@]C�Ęz>m��u�ҝ�>o���-�(���1��o���w�C���-������8g^J�m����i0q�%�[b�T�۰~�*�X�|���)yG��΃��W�\u&k@��Z�Z��4�h@ϲ��eJ�6O��h�+���i	��HWfe��(��`v�HC�"�\�(�I� {["V�>co�^\~��5��/�@�� '���O�Lj�4lw_�L�Qi7������]~�gnLT��,��,zp!jو�g]I�7�"��3�eH~�QL�a��*t{mw�X!������7��)z��������E�6~_�֙�
�W����n5K���	􊔅�iLװ�ZJ�A�����)f?�����K��E>��U4��r:*l���,�K��\�g�J�5���WWo���qb�g����'���5P��E�<�D�r�+����¢(j���=s3n���$o���3F��#��D�1�6-1�|x"LXO�-�N��r
�Xt:�Y�i{�	���Q͙Z�;�f������� ���n�VG��"*\���
���J���M.v��=z~!=�B�K��sg��Guj̀s!Z��L���ǖ�ŋ�g1iFq����5eL��z.7�o���m)a���E�6���wuM�:o?�ܻ/f͖1�����6�Y)$�e&�/Z|cSHp��:�1�RR`d����4r�o��p%�:��ӍE"d�<��Ym���35�2z��.Sxa�|��z}ǹ�W)� ��ң�y �q?�t���𚺟�6���A�6yX`�'~fd#9��40Y��?e'&�§��5�\�8 �����H_w�Ng�,��Hd�)<��LT�#��en�b�`&_H���ܘA�}�"�9��B
l��Q{m�Q]TC�]�z����Z�k�����I��#b�{����`���go��π�ZX� ����� I�t�������pׁ|�^��e���T_::�
���?$C��3���qV������2D�-`��"�����mX�����7J��@�ϔd03�w�t�����I,�3���\}�KS䁙{u.��T9F.�j�&�l�/k~z�!�G���m����?pqoT~y�ȕn��#ٜ�������W ږ(5k�@�^~�r��v��ގ�@�:�^xE HZE�lG�˟ni���C�\���͆#�A�7nh�x
�9K�K�x�	TO��V��$�w��:[T����!�2+U�dh\�W�����Oƭ��s�t�3ݯ�=a,�#������g�b�����(%"��+��Qa�=��f7��j��%��c�q��#Y���@�L�/g�S����Tl�
ݬv�_C8�Ym'�܅^hD���C-���]��a����n'���������6�$e;�W�Ak���{��U4��岁ZS%�|�*��|���@}E.�cӭU|���GiJe�5~�/�,`
�ǪPd&ה�(��z(��j!N.��n��"���?jl�����vp(1�e��+]���(O�ufR�oٺ�ߤOW�m~��:�m�pyŶ��$��