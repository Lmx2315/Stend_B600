XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���:� H9��Jm�q��V� �qc��C�!���L�:[��Wx\Ȧ�PX+��*v���
�?O2=����P�N�8�n�l�ZkCQߊjJ4����Ato@�J�3U� 	G� Hr��c�{���e�mJ�9T����ū�¬�.����u���w�.5r��[X~�����?4j���A�E3����߃���7��@�Β=C�ɫ����VAʏ�S��������n,YBI�n}��d
B7��*�!�sC��<��f���p��z��+wE���4EQ��	7Q�S�YW&�=���|�yU�����M��:;%6�نɇ�H{�.�T�����>��ͫ��)\X��hV���l �ǽE��������F�aoe��'��c����Ǻo�K���"� 1<K�/��*JZ�_�z��m�vR�&��y$�`2�"�r���s%��_�`�ȌI�cwJ!�uo/�]�NYg~���]�Á��l���>�VV�\��J&��cP��r���"�[0D�^�S��ʋ��E�1���	E���|�it�
�5T�`��W:��(���+ @�)D8'�mP��h��`���`��}{�_��gP9ڜa�u�6,S6��XĖ`%{��i)�Jb�ac  i�^4Z�������g��� Ww�����x}0�V�{�������O[ ���Q)Z%\T�Ji�m�v���k_���\5����tsZ�@%���fPWV�mRm�8�XlxVHYEB    1d06     5c0�����kx����2�n�V�Y#�A5d�-��!������j���Q)�����)X�:�x�;���X�b�|�_�����Нa_��IU�QY9N>�D���	cyf�n��_G��T�bW�C�H�����B��a�q�O��Ul}�T�
�E�o}�o2�U]��i��*��98t_�9U}ޖ�k��B��X���EMFs}�gWFH�0��v�=���>����g�B�/.+�:|�]�*�2Fk�FM������՚~A�vw;}�R�}pf���\���Hũ�A�����Wڂ3�F $E���Ʀ�d��2��sl�XBt�o�
�����*��2]%���,��=N`�p��dp"nl���)�ƶH���!)R���A�p�/�F6�\ٺ�Ndʹ|�zi������:Xw�ܛP�90���Z}�Gp\^3Ќ���txs�>�J�혰�m	�Gó�!A�R|t�i���W+ѥ�_7��|���F+��&�҃9�
j�-`� \n�X�]���x���,b�w��ur�H�	숼�Ta�g�kd��Aщ����L�.�@�®������Q��v�3wp�l��Q����y-��Qd�������K��R31�jv�^��Bٚ��X�
��� �d��Tiru���Ry bBF?�4�}�����T+2�6�v(��R�[���߳�/��F~p���/�"���Е��������5;-
GJ�Ѥ�ڕ�Y�w�i��N/�`��08`t;4Άk�w_�6��j�S�݂�U�݅��*]ݒ3y|��N��7��f�
�E�Re?N��:#;>�E��t�����TL���(�ЉE9�&��g2U�@$���v�[�1�!b����N���7�]�$Kq�Y�&�ʚX_W_�3FЫٯ=]{0-��k��i�M�b�		��ix� J~�;5+RR����Ԟ�-�/�g�:;��7�����2G�s����?�V�W��'|�b2H�WE~�*=6Y@6�������_�H9�J$Q�ϣ'��Ix�V+u�PZK����U�y��~�[|�5�����h�p�[�)be�R�����K��.e9:�&\N.�K��`$��FC�L��:�&�!��_�<�gZ�n�5,	Wb�M�� BF��\H�mA�>u����׉2�C[_gt��Y��zW$��P�/�R��۞l0Ѝ6�����L�h� �U�M�|��(�vt��W4��t�H�I�H:!~����1Y*�b�Q;P����a�j����2�Dbޞ?o�)��J�+d6��/�@R:*����`6�P���L��;��9�c��b�I�C���S҉L��-�׼1�j�Ez\Gq��B\�?���6��Z�k����l�T{9+x���0��M��H�N��T�Pf+�����c�ʼ>��ϯ��J�]D~��R���aF����|^z�D����O