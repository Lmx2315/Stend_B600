XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����'+��y���@�j��H��VGơ	AA�i:�>Y�{{�܎�8��`�-���ݩ�`>g��BI�^���"Z�aQ*�S��~^ro[��q�U�>��4�2Q9��`IDB����^p,ڊ�0�=���~�S��u������*3��)2���q-G�L���;nc�M�<��ԚH�D���O���~q�V4��&.�X��M��e���ͪP���*�Y�T� ��O�B�G�(�w��ޘXU�y�B�������N!l���9tjt������<��'�EEu0�)��ճ�	~{d�È;�&m�X���"��o��n��K�m����xQA�#����v
�����<�'�Z�|�
VQ�ei ژ�W��q�:��˩���(�H�1��@V��_�M���}�O]��
ꐏ�5�k�D����/M�Dޫ4��_Nt����1�#�����a��̲$����'ؤ��_g�K�������~�i�;%�wzH���ڼig\�����3�_Q�����ϩ��1Q�B�Q51o�,�ƶ���V��Y�\��������Wb���׀�-4	�7�G�	,)İ�|�m����ɼ� ��]W�nېN>�C�zb��W�*9SxmV͋�*lm���,�8~j����1gXV}OT��ӓ��^2������u0�'�a���oJl�H���5r�\��#�}܏v)��w��F��g���B����}3�s%��AR���d@-OX-���ݭ�h�,��pr�jWОt��XlxVHYEB    1001     490J�'P�@�x�����S9'0:�,&sp���Z�J�փ�U�Gy>m�G��
��$�A0�qܘF��o�v)	�&�`,�b`��t&<k�� ��w�0Z_#�jCT�e��VD]�LL(1�6 ͊Z�\~
^������3)�)���}	a�^�ۚ�a�!G���Ǎ�dl��4׻�MEГk��c���������e���$w��j�߃��G�Z���k�N��a�`a�,�o���0��0���H��~u�.S�9.楽X��S�v#���q�[��if�g?���b��pr��z�d=��Uᓊ��ru�����=p-��$��D��-��Wޝ܌�0p��XK�]t�1�1�!E=��D�r0����<"������>�2�[F�XqIE%�$
z��j̧�4x�(����i��,��/;�J��2	s�h5؃�ҳ(��f��ph��\�?��2���sY��-/4d��6��#��{����o�S�&nP��Z��I�����_� ��fڗ+g�zBΠo�j^�r��J���f��q��(6ಒ�C"e�ƺ�E��ç
�di����Z�Z��g~q9��e�o�Fv�(&�Dx���{4��4m����#�ܚ�9�[�ڒ��"�-�o'�p�dV��]������RUeH��ذ���6��@3t����(�v�*W疺X���Y��$ �W���MgG�J��֊�wO��qq�U�ܮ	j���NY��~�m[VS�rz�j�l�M8�b~A���T#�
���d��|�``����)$���!@�6�>$"@Mʹ��~��KEs`�}\�3(jVc{*�!t��Yw���F���b�W ���MsB@�Z�����#k^�e�S�el�Yxz�R�,��F�8R˔X�{ӕ���e[��ױr��La����I�d��D�9w�3�N������,.B�%�W�5�D/�����lMt��"�T=�j}lK�f�z6ڮ$� �&'�2l�G��ج�/�Ԉ��=>���Y��!_e��E�2����W�Q��(/��=J�V��h����v���(�6YO7yR����kZĚ��!N�<ٜ�. �T�����)��q�"��S�`{�^�$�-�ir���<Vꎙ`�I�MxJ�ʀ����������m� ����