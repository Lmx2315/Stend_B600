XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��͡I�h��
NTW�Ё��i#����"�]��?��#.��/l?S�.�E6�Q��jŲ<Eb}�y�죹,�{���
+L�mܜ�@��<l�͗�T`b\��m�p����'`�Z����(���(QBj�15qg��w���;j�l���"��±�@����E��G�`�%��j�0:�"P�����+.}V1G���6��3O� �I54p�w���aZ�,E�I��<7rQ��k^LNc�낮`��B1nk�>MwȚ�&�D�$2M�[��2��4�TN{q���b���$`�����2��C��קVf%"N���Sp��w�i��$��@6h9H�p�Qff��-�A6�[�nD�ͥ*�d���Vj�~܏������s��~̼��Z�@퓚�:�p]Q�lU�5abNY�m��	q�C9;ң�`uu3��/��yd2�%b|��^~�kt�*��o��&���m}w��H�v�Y��_�GZ5�9��jN�#�A���wo��@��&�Cv�c��k���Y�����<.�hT��Zd���0�#��+ "�i򀬣z=d9����]HH��^���7��ygf�<����%��c5��"��!a�j��$�1��⫚>�6��˼�`.�!G��m���� �%Vq����}�J��q��*`��B����=!d���b�p)ڿ!�M����� .����N�)�Te� ��Vq�0��;���8��.�k �,r�������.&�o�#`5��2^J�Ƚ��jk0��X~
o�_AXlxVHYEB    26e0     820�#��%��%>���i^��]=�j��l�0�B��n.�f�yX��|��;���r� ����ǥ��H���,R�;?l:nx`���R��.羦b �s�����Δ,R��.��o��RÅ�>Z
d� #e�\�Q�<N�}� ,+h�&%NVr�p��bc��������$љ����� �t��A1d�A�E_��K�� ��h���n���N��N���2V�����4�Ő�*�r�k`�ÆOs�@=`�1Pf)�ND���5XM��4F>���02�39�1�%�a�<g{J�;�E�-�(�����V��l57v��x.Zsf�ϵ�m�ɚ�f�� �����YH�b�:~��ʎ��z�v	���[����b�|v��\\D�*��_#�5�ʎ�������Ĝ �T���6�\$t�x�5J���P���6X@��~%��#g�]=���Pg|weTeB��YOm����
�s�e�C/���F��/�������4l�Opa�Y�4�T>�f5���.Z��7Zk8������+i�����'T���+z_q̥P�:�al5���r� �%���������#�����T��[�N��lA�ˀ�)��T���i��WF�n���N�*�3���m	3^vp�蹤R��ݺ%�0��� �p���`v�NM�C'U`���̀;�Q�Ȥ�+M�SN�LeQ�0fܞUVMFCK���O� ��߳�P�E���/�:�o�e��"u��?]9�#N>�k������e�+�@��F�#�>�E�r���o�x9������}<��i�q�����~���i�u!�t��A_W?(��1b�i4{:f�`����gf��%�evW��i1?pW��2Y�nPm�w����Xw|�٤��%OЕ�f4E�~���n����5�9I
�6�d�����FNU'+�]���s����)���Đ�
����鴐iEvB�"������M?�e><�[�Բ��S�ڄ�mV��X��}1�ȖM��̨o��ݟ���(ՠ.N��t�e�uA&2W'l-\�w v}f�O�����Q�Y_��̜p�G`�GN/9����p�I6hL3�
}����� �"�+���F�p�8׊�d}��)��������`K$�7�С;K^��$�7��|z�%F<����e%N��IrJ뫚����z��rz3�~�ҳZ����tH��y��+�3¯t	�7��:��q��B�o�n��c���vfT�x�A����cz�0'�s��@0�Y�ޅ����P���Ov��z��Ѳs��X���O�qIK���t������04C��P���ۊ�{0�4�Uy��<������|ɚ��5w6��_��S���l���l\��v.a;j9S< ဲ�e4�1�;~���Yk���C�����JY�P���[����D�3�4rR���X'�x��.dy��:���n�壜�������r`�̡"a�'�]~a{���uOP�G��#�ێ��(i
��?G��!5]�Q�`G�8z�c��Jh���^�~-m3���뙊?��y���k�C^�+�~�4gc�eܿ^�	c�j�i����=��q����݇�O9�"h�^�9��1�5�۳�O��)m��Z�����ZzZ���̳[��}������e�Kp��o�۝��G�S�n!����.G!�֊��3X�dĺ+��4�la%F4�Zɮ�|��b�ϰ_�wf��sRK~H�]w�بQ���t H�K�����^�j��9��� �~+k�vYlB���U�a���#D�
ڬ�$;Fa^�7EJ�1�$ϗ=�%1�U�G���%ą3�u1�DZ�A�>!�w�P0_	u�"�̕�>5���"�P���Ͼ�8E���@Ndse�=x����� (�v�Fl�����5I/�Kwk>�*��sLA�l�U��0��M�"֯B��J�����!׮'=�^_}rOW��RY��6���ˣs�4Q�/Np �2/��#֛��?e-=����a�7�ty�6B��qfF 4�@��<e�z�<�K��|�P编����B��З<A�,�U/ 