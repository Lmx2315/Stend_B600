XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������&����"�IB3�r����X�)Ϙ���o��kt�~爏M�&dUm�;D�\���P���EP�T?�X�E+�<W��4I�X{v�<�1���!;F- ��H�/ ���Rע�}@��2�j������_��b|=+)�6��(H�8У�rʺ��^��zS���7.�`�Z�B&��V)��M���q���J�F���O5k�|@lf��8��)G=�`;*@)��f̄m�6���h�_KE����v*�;b�B7@�o~�Qi.��*1�)l�+G�U�`|9�!VS3a[���v�k?y?*���dԮɲ���*1�Ǐ��7�>а.�*��hf���`�L$�=��8��8��{K����CV�,H�K���=n��$�w�����bG�?��og�9�=���M������}5m��R�vR)���0�︻K���z!���W�{�I瘇�ϐ!z��b��D���-�ҽmu�n+����P��aɍ�g�7�6�% ���P}-���� q�鳐붘���ܭv���/�=��Y,z����(QA�.���x���!`)E�Wq�G����^�z�w�$!bB�.�7Bv�����3;�G	B%�����{HO���B�l����*���C�������l� cI�����'����N�PH���A����)#y�m�4c�0�e�����[��ZjT�V�C�ɲ�K�C���� �s�	pD:9C?a�:�}���XlxVHYEB    1041     4a0Y��Jx'\+т4j�z�����m�8r~j�6���1[S��N������@``�[A�!�CQh�y��}�z.�<�Jca/���\�)���5�Ȏ�8�l���3L/_����\@��>&�L��9T�t��ō��$���48=���w�K%�KcYl>|s@V�R&�ϕ7d`_���G���F��R3��\%�bi�V��f�#�^}�
���o��t�A.�]��i��>D\�-Qv��(���n��n
�����]E-� ��
x#��O��&^VA4L���v�bWƒ��Fɳ�B�XvAsB�x^鵫	%�^�)����J4�̶qW��\��[�n�&l��x0���q��>��rc�P�t&��9<���bea��OùE]О��������a˽B�ʬlBo�WQ�殾�*��%���.�i������團uexS0�����UI�6��!o�>��wh	]l ���yl�de|���ߝ΄��gĸ̌�ѭ���� ɹ1ѦmY�0�A�J4����SOb�X<�y� dA���G�.��5�F �Ɋr���\�z8`�Z�T��9f�r	j��\�G�{z�3�����ɃQ��^.|0�M��7�������1���4�b�\���t/)�N?���p��&/{o4�O߫\�����b�.a�ը`#lN6L>�7��ۀ�w��P�CI��g♓NP�n�Іp��W2�R�e'��k�>(8Agx׆��HU�X�ك!;B�rK���P��z����3��@ (����&�����̽�#o���U�s��Fewn���?ך��ԒQiw'p�1��cL��*&t�d�l�p�"D±�Gu�ܗ�A�jr��g�����G&4�$��/S��	̰=I��b�5#1l��*�8�9x���+���X�iҷ�WD5y��'eubg+��K��O�!�a�� _��=ӈ�ٔ�0h�F���V�|�����M'�Zx�	�6!��� ������-��|��J�m �l������4�u%�N��ɛ�lB����YK��1E�����
�n��,�l�0P�l�UT������
�9s|���.�F:]�ج���|U�S��[d���6�~I�ox.^3�A4��cS}���I�7�[�{�]�0�������z��������� ������C�>�3G��e%���