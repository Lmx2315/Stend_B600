XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���`Fl���eU��F,8�]�Z�
&.:c�f��坄B�Xcb�yU��a�� xh�d V��������d�*��� 1<���(����
�(���tN��nh^�j��Ǘ;&���66s�$��֭&ʵb�)�T�x=��޽N>�w����β�3C8�Q��bs����yG���s������$3^���(f�$�"���.��u�.���G���Z ��|����n�6���?O��\��w[#��lA}q *!vQ*���K��a�W0��I:�Ip�C�K�]��׬9��]��d/GS��m�[��{��e��4�����Z���Ț�\�v��P��i+<y�؀?�I����sB1&Fץs%��s�  �H�stҀ��b[�|�q��k�$3���w�lB%��������Z�罤��8�[E�%DDI��� �T�:H�'trX��5��@�\o*x0�|0!��qz�U�k]�A����{q��HZaKK��n~V �q�:�]qpW�<_V����]�,������j�<�\�&��� �&��G��fH4���:�6b#���,�S�J��q������,|vN�}Ȥ�D�hVA#`�|Q���h͓�� ����+� A�t_30��0j-#F� ��kz�p>�Zf�2j���7��(1�)@�U�m��'Si�n� 6Ր.�n���KV�X7 ~��!Z�ހ�f�����<<��c��;
�/g֋�������}?�Tܪ����t#XlxVHYEB    152e     580��e��q��U��:?�~n�Y���iq���D��!�L)����@�8\hD�#�C������I�\M��,�`�5�Vg��d��ִkW���3�%�X���� e��Iv���ph}�
si���MȜ��r	yk��p3����XBL���>���Kwq��^�r�<fE�O�K��K�B~G��P��n�r�=^�8�M�0�A��BT��e�n+�wW:����yG������y�U4G��c�ut�\�viW0=��?�3���)�?��V�1CK-�g�M���A ɐKņi$ݲM�,-��>N��G	�D/	꽾��ߌ�@����j���q�'%B�8!j�b���	�Jq��Q�����3޾��[ k����e8O�)���|0�X���C�@�����?�#�����P�[;�[����`�㟬�Et���Tˈ!�Պ̜G�5c���ࠡⷥa(���:��K�HM�j�5y\��Zng~���ΰ�/�hrl������xzJ�	k���H-�aqҍ6��#���W�
�h���P%p�"����9�����x{�t�#�Q{�~��$�c�5�U�oP�5�<�-#��b(	zW]ND���6�D�����,I�ۛ0���$�#g��?r��ٗb��s�/��G�'0a.ԥٽ�N�4�.�;G���K��п�ߣ���̋aȺg@jngv�1�n�|�a,�X6 �+�
��`r�Ǩ��bd��y�:� a�JnV���>@XzԬ��F�������6T����Hi~��"�I�'�m�>U*[�q�1��J�uL ׄ
�,Yd�k΃����I�7�E����.X{p��,�b��'8�p��N����#*to��U��$�y��Zc!sW3J凖Ti�j��	5o�6}�M��=ͻG/��o�~'3������̽��?C&#� )�3�3�+�������z�X�.������WĲQ(�*��u�#�sW���FP����m1}N5��n��@��>0�[��3�Y��D�R^}�$<7Zu��_���wS���L8N ;<Ρ�������j���0#��XDGR�|t����K*0��@vzS{H'�7}�C S���|N|�voo��(C�I�4s��N2��o��?���m>���d��\�p^4-\���0��c�\�$|fȲ*�7�����լ�)l�b����̠f�>��N
�)铽�++a���[��|����m���k�mEx���JWHg���!��	.��!YXR���7��<��C�5�*�K���O���i��(GfUzu��%g�/���7H�C�{��y�g!��N���O:���qg?VG��A��0N���6T^��,'蜑Xiީ6Q/f2�W