XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Y����w@$��C��Pb���	F}ݲ0�(7P�;��sY����($�t�(zMq/���,�T*�4�����a��vC����
�r;��`` }�i��K��@9�؋��U�$�4|�&>�����8v�(����(ݛ��艹���+�Al�z!��	�7��p�,���@'�)��7�8��n�dUv4w�O�u�� R�Qz��ft\�|���u\C��;��[���m�
R�@fo��H�H=]�k�K�J�M'�qMu����xw�2�X)����������"=\E0-�'K�N��G�8�c���a�Sg�f,(Q��4æ,���͋�N�@��M����E�h�~���@��;�2�voR��4�p풄�Q��Z���΃G0�^��w�ӁeΨN�sGV����̌nS�W�X�<��j�+qqP��2�;�M ���n}(��K�"ʃ���z?-��°v��m[%�ЦE��=x�t�,�xYK�?�a����M�"�}HJ�i��;%���ĶZ,n%�-�\�4��n�;�u��#��FI��I�D����?�\�&�p~��jN�����>��,��a�����rj�ߠ'��{xҲYS2���/��ܿ���6�R��y��o ΣЂf�6�4��	�!���S�*�>�V��~�d��k�ތ��� >�̬܋A���Kg?FNda��;���U��P����\��˃ �5!k w�:�rt_���N�"�Ih���E��۩��}3�XlxVHYEB    1902     730't<�#r��\��aN���������d%I��c��Pn��(h��D~Ll�Y8a�I���H��j�4UW�R��ī��U�����L1�l�:~
Zo��:G��G+{�K���R��2a��L��8�$JL'���.{$�z�8M�L�9�G`��%I�\l�};9+Q�f>�#1�D9�oy+|y,��c���vz�wKK׾돎��m?S�a�Xk����x�ge�����\D�l��+���f�C����8�iAJʴ�)���CTktW?Т�G�4��y݅��U.0i����"�6n�cy�H5�Z샆�6L���Q�ݥt�IkZQaU�\�%�?�k|�2������%�q�/>��К�H�Ah�i������* R��&\�TS�s*�37jyɠ�x�X�[�+�c�������w�4��z��*�vt#\��i��X���T����8E������! ���蛔��»�f�:T�1]~(1I�R���. z�]����.\�z���|b`z��A+��F�G��p�p<Y�fSǱ�2hR��74�-���[�:6WyQ'���\������ ���o���ζ�����,��l��8I����R�bvOmY�(�	B�1�q���)�51��k�Z�kʓ'��/��`�%����s2��6�gz�{��	�L�%%Q;�����6Klx!̩(�lErH��=�W[��!W]��`nk��f4G���}
�Ǧ�a;��9 ��,������Ӥ�]m��%ZA ���V���$�G��^�O|�oQj� )S��|X2B򠌭��U���U��	��T��)5�k���l�.����:
pf�$����Za+2	�$a�qg��B�<X+��� pF����ŗt�,Mhv:1eZ|T��R�r�����R�\�A��U.��̹j���r���`�������21G8x��{���-N����g�:VaP)5L�L��Xǈ�� �v��H,<E��*�D�gpFߣgk=ӕQ�<��o�,3ߋ)׎S�9o`�	�Y���o�vH�~!�v�/%��u���밟k;�d
�7���p��*�J��7.���׏(�WN+��T���Ǣ�\.(�x���M��$tt~qG>Xy�	���f�~�9Hζ�%��(Yq�%i��	�Ld��&�D=B
��(}�th�~F�'��*�޹43����r۩�I�~�J.�m��y��H:�y�M�u�(�ݧ\q�$b%Z"�昴D����3�K$oo��(S��&
eZ��`7$Ѷ��Б���[�Ydd�)�aL��Wn��K'��
�qQ�iqe�#q�7�5ԌS#�{����Dk^�n�O�*y��o��>���Q0��g���\�6X���q�8�B��c����^v6,3S��<�T���&a',�9��xκİ�2�����`���E^y���c��@͉� ���&�}��Q^}�����\�^����&w8794FuH�d:ō�T��4���٧1�P@�Q�䥢�E���o�Y��ƥ�U�^y��`JЂ���(;�ؤ�;�%R�y���Xxz�Õ��g}�v�"����~0��{�>�����5��W~e�B�G��1)�)^�Y�����<�r0x� �� V��F5A�e�gVX�ٯ��WT��m:m����4y��pY����3؆�䪺����_^�����r�OIy�]Ŋ1��Ӽ�r?��A�H����mK�w,9���/}߉'�&&i��IA Q��iC?\r_QE�X�Z.�Lg���l�Co�l�ѩ %�<($���d�&'����C!K* ��