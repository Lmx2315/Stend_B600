XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��.��`p�0?�
+4������$����0)V.�v�&��`�jD����m�m]>\�)� ���wp�T�9��>��ܣC_��̽+xR����¦q�WԬB�(�3�-&$�.���E3�G_o>
�e/�悝�V��ԄF�ű]jJ�:}/k^%� �p���P�J�}�>+Ma�b�7�oe���C�!0:dϥ�4/��L
�_��qQ�T�[| ���g�\4���Z'7�Џ���d�B���W���dH@��$So?Jg�/�Zn�-�`��y�i����Z.�r���3�(��sr��ۄqO�xߛ�:ĭ����u�	YO�N�u3E�ߒϸb�_P~�qt�)��	��O��n�4	�o�׮���������d�X�hK� �\��O��8(&�'̝�{!&���� �� �k�+%���0��ZԖNan�m��n_�_%T�"ȳ�avDcZ5���}�%�e9u�J˚����"��@`S�㾸F�ѬL,s�����"w�t�껧��O3D,�6�Qo+Ƽ��O_t`��0�o�� �A�b�|	,�S�o�t{7Ap۽x�T�8�KK�V�h�3)��8у3��҂)!�/�3�<�S���+�)X:���*o��h6�B���*D�[����0���5�<I֩G	�F����Ψ�Oc?#���V��&ϕ��a3�U�s$qe-6�8v�Hn��MA�C��N�4G����'��=�&8V���M��%�xb��8`�|Vf���%y7��s��uXlxVHYEB    41a2     c20�؂��p�W��* P�����C̾T�Q����n˘g��v��h��!�`f����DB@.�81��g~%vC���p�8�������!��L�D� �����JDA
�������a���G�iF#���dU�yb�H��u����	�m]fr6�����>���|����O�p2��N�#W��*oԷ�P����Tm2�;��n�I���ͤǜ�<v�/���q2���ܜФ/~f��3�ۣy���#S!ϕPN�)t��]c�X��rl�F�Ki��!���R���[�ߢS���<��W%���\����E�S��&%*�
!/��'b��ol<,�̉��[�(�{�V���Rq�>���W<f�.�|��TޘT�W��-r�v� �	Z�.K���XF�;��� �A�cr��|�6
��q+��tO�X�"�-�@o�渐�.;��hD�\Vmh�VƆ���{�\_��m���!kH�@�J?�F�l��	��E��̄�N]o�9�	 u���A�K|�0��ʤ��$<VX�����!���c2~�G䤡�)'�M�I�0o\�-��u�t`�e~jC�aL�����&�lǇ���)g��v1K$�����ZLrc�<�8_͗7E�S^�%Qaӳ(h�oҫ�9`ܹ������2�(�u�Z�pp��l�!y��C�Mv��gq[Z�a�Cq�pGt}@��r6��@�/m�v�0�Z(�Km�?E�%���п�3�����:�t�X2Lw�ٚ��LG���y�%^Y?f�Pm����d"S����n��`\e����~G[vl���B����s_�{��]��a4�r���AX�Q����475��ˆtm�����$6]�Zp=̰e��@�F��/��Ld��Jv*Y%w������ʛQ2��J���8寗.}3�"��͢8�/�����^zA�P��%����mЇ���uI����@�n�<M��r������{}���?"�~~��5���,��TM+W��ۭ��,�4I�����_�"��Aˌ�d�蕘���߁.��צ���ř;�(��׏;V8����5�E��Df��=[�����ؐ{�gc.`�?q�X/7�?l0�l.����;��0ĀU�M?�k����9���+�zQGt�����IK�a�̬�9m݌�ƾC:٣|��~<n��kp�1guOE����޾!���6+����m�-��?̀�H�D$Ӊ��#����P[G<~�[
��R���ۊ��΅-���p^�?���w�m0@*1�T��ߠ
�Ķ��]cZ	w%*A��<��ȕ��>L���E����I��1�b�]2gt����y�7L����g���z��N�߼9���,)(�`nLS�u�M��jL��AA#&K�-3�A�1|�/�]	���[�h�ň�l70&Q�C�*�?_J��Z<�7�$������9�KoVY���sV~��;��5&(��]��9\�m�:r�ƌwQ�|!o?��'U�g���T��~�mB��r����<��L��5clv{&����j�. ��T�r�n�^�$�#�x����Tz�Q�����ਧ�����{q^Gͺ��ڨ}�9٧�4aV?�\t
�i�5�>���R��@Ks�"���Mڸ=�b�1{�X��P�2(%��ڎC���~�]��lȎ�A�Z�N��mU4<��DA�eLTM��\���}05r�PS�Ȅ,s�l�����q<i�9���b�ׁ�|t���ؚ.B��mʠ���|����6����[�;Pi_�W'���$TZ�dZ�!A�U��k	A�I;���x��ٱ2ON���w|Jv&21E�آ��!��,؞v.ţmq�c�z��a30��З�Ss��|��)�G�σA�X'�������yf�����Ѷ ���x'�"]9��I�����AⳬaD��}��?R�e���@�����Ez�����}�%�cv�,�gs�HjY�1,�(N�Q��o#ր+�O)w��-�q�C4:��[9�w�tzg���CV����� �=��92ޜ�C��SsM,V��1Ydh<a������K�������7K��99W:7}���Ѝ���l)� Gq+a����ȏ�%�:6��K8�hƀ�]���@�%gHuu�DV4�2K�ā��Xn��0��jp�&��OV���?���Е#�6!Ҋ�־���©ʥ�*$��8�xG )��d�ݔ0��4��*z;"��A�c�,O/�eou;����8|ڸ��$�IV��I^����[~��K���	CeZ�'��fNSG��h �R����"Qt>6����,�P��!�I�0ʍ��d�Tt�ĆR(��JTP�q	�Tq�XV[�;�[���<�U����`��َ�_��v��Mб;H��5�p}
��vNv/̘�͎Og_C�%)7��C���o��m�� �o&����rx6��r�co;��
q$@ˉ��;W��0��G���{��8��UU��9�zI�u�T����F������:�������qe��nI5��`�wt]���mr�N�+d'�RNhI�4;ǟ����������yjA1Ή���^�ڧ�b{��S3F�prN%��}��LNu�5��t�Y|����SaP0����j� ��
�0,y.���΢�P(��V�w�{����R'��R1 ���$��
t���I{�*N5�\�����p#>3�� � C$��ff�杯Zw�覉�,��-�5D)�DP�`P�ʨ�X����+�p�!y�v���D�".1��Y+����N}T"�ђlz��+SCލN.�X���sj|�U��ڜU��OV�U�Eۼ��Z;#��|������Ee4�z�|�z�O�P��i8�Z^�ȐWa,C������6{´�B�ṡ5
���>f-�³ �˜a��#�l�ʝ��Q���G�V
t��Xi���+O��YBߏ��Xq�֦ms�\�*�8�"�c�[�I_K��3Ӷ0���2��Gp����Z}�u�o:������y5dR �K�^ P
G�e2n؝�}K�