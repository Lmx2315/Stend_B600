XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��\�Ԡ��4���SG��D��/#P�`i��a����l� ��+�0�HQ��=H5�� ��E	����E�H`h�'�%��ˌ���
�K~;P���s	/��C&/v�6���I�G�l�^�4���,�o�	��O���6�����}'��7_��u��@x9��m��K9�Q�y���E%^p]L��� k#�ҍ�A���������h�B�H��$T�+l�P%�A�]S�X�u�a�+JZ���yTI��U�$h%��l0:�I0)6���	=����^$��$D��/���΂y���k1dR���}��EWe'�g�����O�"XL�2�{��v`���(���ʖ�.����^��-�cS��]g��� MCd≚����vWs��q�y]���M l��>���=�RTV� ���uJMŞ�$��i4�k��:8S��zMbhJ���{O�U�~&�f�/�`�ݾ�I���d�@�48F��jj��?��
�G!�,��jS�)�����+�R��Q\�/9�T�|�g����nc�L@�H������f7�W��u���2�}\|�P��q2�c#�f)�r�|f�m��Ex�8?-J�Զ�*�2�wZ���"eO*���ު/�A�V!T�\W�>UDP��q����S@׋X��-u-�8�we����}�%|�x�G��W~��Sjׯi�o���i������/{*�}i*���������g��JUC ;��p��Qy���X��zqSZ
�[n�M��<!ٯXlxVHYEB    10ff     490�H��{��<yl�f�h�o��L���Z�-m]I��j�O���b��Ɣ(�g���j~|

�]��xm��� �&D ��+��h��� a����h��h�|�ĭ�2N�F�������� ��P��rY���;��1��S� ��2�h^|���`�����f��I'*���vm~N��AP��v[�
BDvT��P/��i�My��+~�G`�U��q�x�'�B���~r�~챴�k��u��5�ql��}ĉ䄵"��b5.b�9�;��4"۟  ��E;�6}�Z��>�B@G�I+Kn�u���Xp��&��4�nڬa���U��#���S����x��v�^N���6�e�6a{��}���zZ yI �`s��ǜ��v�~`��<���/Ƣ#/���Tz�
���J )��(TG2�op����P5�&�rx��Ӈ�њǥ��.�񥒁���fR��XV(W�Z�]-�H�o��JqPE��G�X~���&�ֵ�R<�ev)���&������7��r��DT�{��XŖ��;��Vt�pf8�N?1ZS� \��K"âh��:%��9��w�@ce,�����o�$����xt�Jݕ𵏥~���z������s��x�
��sYg��dS���S���N�|ꛀ���O<zJ
XeGG!��tr�,��4� ��JֿL�=�C�=8v<�g9��-�`�	����	�[�l�4?��gvn���B{�d\CN��i��<�-#��kҌ�KZ������n�րO_q(��ln�Xl1��5�P�nr�Z�������]Kq��!�M��*>�C)�.J����jͼEV���G�q�)�"7}�`�%)*���*X��ʱt+S��z�|r��_���}�M��^�BB=���<{wZ�ț�f�����|9*mx$xE	���!������t�E�%M������P<�z?��_�k�R�#I%��vPǨ��Ѡ�אe="���|dú�d"N{��W�%�d�y.�;�����|p"�k���v�|�>@h�sD�W =�b��?�V��N��5L���*�_6:cM]��mRP&¼�!>Z	�Yd�(�{�&$��1������r�	���+]䯵	�����/BzS!��:m/N7	�j?��'�I��6b��iz%m� ��k��&o�k�