XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����3f�D5�i"�5��Y��	lƱ��<�}�M�Q�b�vJ�;&�ރ��Eh_Z���֌@�Vo�b4{�9���Gb���;F�1~�r�,���G�L�_	���(T�ò��8�����ܡi���&�z�v^��#X�=dK!��h�Eۚ���i;iܺ�!U��b`N�+��?�\]S���~@�9����kZ��i���ާ�#El�y��3�?���E�p��N����fR�������P�K��z.�����M�:�̺3*҃|q�Hu�&����9�x:����N����v��8#�n�A����냕X#ǥV�{�;s�7��@��|�R�ؠ�5�z���2�� �c}��и���DA��wvf��р�9-θ�9��o��Y�'�}�\Ũ��P���'�&�Z�|(V���T�݇�L /E�^-���������n6�nQٸFܐ���q}턭�h�H�,����n�4O�%�A�{r���vq!�*1�D�j�qvɣq�P	���cT ��1��|$<Q��6�������S�l�ul��O$�ϧ�DT�*L��Zm-[��!-��3V�;�ur�7�*Hw!qP��������W��(WBG��U�Ï��O����O�D�Gv����W1v��CZ��5�x_$�X?�CY�p�\)꧗mg�	��R�$2�k�E��@����+�rOJR�/ɸjîQmb�:�ʎ�G�}�	N��Là��t��Y`�p�⃎1a�w�w�/qh�nXlxVHYEB    458d     8b0�v,����g@��-e��(Yٍ|ˁ�B�[�a��ښH��:Ι���~8�����Â�Q���}�B}C��>E��
�/Ǖ���O������č3�Z�̳_F�h'd�M��܌Ȫ!�0t\ׁ`�an'R��53T�U��I3K��֔ŋ��9ʊ�����a��Y��T��1'J�����M�e�P��V��4�CT�E�*m~��������5y����d���id����/���'�"�L��#m~ЖG������
�� ��!�CKp;3,_����Jto^��rK*����=��گ`�pn|�u��v�ﴬ:d2�(���p��ڐ�ւ!~�K?�\��hs�O�"��nG�S"����S�Y������9.�
yP��%�5^��/_�'`֜���6����;���@> �S�]�¸����.� ��@���E��ب|��ӈ��l�yN��G�8�z�����e�*n{��x&����K�A����Y����4�hD�YJ	R�$���fv4�����}�L�}/j�����HX��"��,�	Q���B!c8��<.'<X�q�@���e((W���t����;$f�g(���y��d��ٕD�����I;{�����"���BG�8$M����z�w��I9�[�k+�Ӥ0���5���»)�Q�dOfrw�ɴ[A�B��DU�; �>!e?��� �^D)��.0O���97������,�3�v��D�8rgu0| ������Ώ��c���s8
��������Z�=4�o$�V,`�� & ���E���u�����F�g$�"�
ֳr����Ѯ3�LJK9k}���}�SA�8�[�*nYXP������4Hn�.�? ���X�}�зn�X針��룰.i�����`ɥ��DtGa4V5~x\/6Ҷ|UvNXg�kDz�������g�R>��M����+QȾK�Q�T@k�b�ߓ�hJ�YС�
l4��}M�y��Cx*�{5���B̼�sf�m���ԕK'�b��	ǂ<���S�9��!J�����cqUB��x��2����k�
�#��%�Qp��y�$����R�m��(��*����k�e�RL��Q���^tŦ����o�C#^XK�ҡ8�g�F����W$Մ"��"���_]����@�h���2�:i�\�]b롑��!:.Ix<̴g��W>B�O�6�}Z�f��7����Xz�����p@�X��@Ge�P�L8۝K�HG}%kUr�5�N�"�$+$_��uA�B۬��Z�5լ��_k�1��� �'�"��7�a��z-��Ռ�+��������W(���}0���۩٪�D"M�ȝ��I��-iV+,�gu��z���e�-�e<Cw�ח�hڿ[g�ض�Y@Ϟ��2i�?n�M �ų���g3N��hx(��B$DOb�vӴY�q����K,,"Jy�2�+�.����Q�_H~�B������/W(H��L��׷�,�9� ���l�8:�~F�6!��_�q�p�7�7Kzp�(�*��E7Ƌ/�ݾ��&��d���j�n�=`7d���f|z{��I��m��&y�����k��m������6u�
�6W�@]��\�:y!��Q�C��Y�R�U����ԝf�>о)�(� + ��j������F"�4������3v��.�T�cS�Z�q���]�6�_{��9P��R	����B�����Lt�K��Uk��J����J)���}�y�d�D��Bg"�:��2m���ʪy�|���8�l,�﯌=����D�t��sNpTq��W���3W���nf�Jʲ¨�X��6>1J.���F�Ձ�<�R6�SR��D����p#��\v�O�ѧ�x��\���B���S��vsJ�~��Y�}�p��/2��#��%�_�"���	zs�%P9C�w����`�Ws}=������CanK�j5���P3E��
|Ȥ�I��PO2C���B�IӍ{XH.�%��C�bb��o���*i�����ޜ<h��`�����gr�+;�4�
��T1�in��ʖO�50%����PL����#��V6~�����a�Izq�R6��S��r���K��3�-!��i�f�"�ɚR����0@�7�)rWMǁ�Y�h�|�F�y� �\v��V�"�Z�c1���5�T