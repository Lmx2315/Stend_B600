XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ԖLݕ���$��-�\]��t���`"(�8�3A�N`��c��z!5���y��ŬX8��pF��@�#ɸd���"�)WGa�ɳ�l"�R�|c�*�����)�������
��Q�ލlz��ç��	#I�Z1�nJifL��:}1���Ľ[�v@P���~Ec*ٛR�kj'�L�u��3��jHh����K����6���R��0��K:�/��7t-�2N����G(��w�=�ĩ����r�8�ƅ�����;��O��l�$�Y��%d����.����(q�2��W�%SVcaHn����h+�BI��D�T0��[���O���u�f�֨��=�)}���6�7�v�x��l�I�)�c�w�k�H���;`�?C'+�iŀf�����D/i~�u�Q��y+��@�]�D:��L\��[�b��:�:=8?�#%��Ù�z�R��J(���bąi��Ö
�`
j.s`}@�M������{E����,fX�1tu� �ʷ��C;ր˻���[Ϋ>���e��Z%u���hz
ٙXZc ���V�e�$Ҏ�8�:O�;�X���z zc}�o����^u\$e]Vi�Ը���}F�.Yⱡp��Є�Xc�!4��~,����"�Z��DC��vA��ݚ�z׉�S�+0�N2���Z����A�Kz�?�2�qt&�R�S>��r}�I�t�,tv�-�Ε�5�wp��� �	g�*�u��Q)�£�%H�(�^�_U�S��"XlxVHYEB    2695     680x��|�c�Zon)��*��B���(��)kK���6e��fąDQ.�c����^�*��Q�f���{@����.@+�&����Ew�\B��OP��Ӿ����A��m`�_U�S|.�t��GP�W>ұ��q�o�j̤��ށq�e�?%�=+r�D�#�O��}��,��\I�)N"��U���W!�S��݃d�2�[k=���=�nom�TiM�C\�* ��$��̴&-�پ>w��D��s�PxA��E���!���%}X���Kz��΅1��t�n��/��"ov7(؅a)��m��p͞�hl,Y��&l��< �o^f��7*֬�w�|(k����Kw���)r��d;7^�dF�>4 -4|�{�5k�QgR����e7�48��ߢ+	�2���{9���ÙYf��������v����^ֱKj+{�Di��Б�~��Ӡ��6�|�=�t�j��W��N;Ħ�J���qI�c����U�C�4�k���jw���a�C]��~����ݜ��=�w�G��=����(�D*������2������7PF=t�~[���(=p쯬&���px!��K���/������X��I08�p헷���Z����t��5�-�ƝU�F��<�_��0M��N��e,#�V��'Sj5[x�u��X,p%d�-.I1�e>R��1z�1�z?d��>v��Oj�O�E�Q3�k�(���`/uǤ��w��2��K�.��JtD�}ϓ0�X֐�*`�y�t�@�,�/Hu���ʘ����H��T�.�9���\�'�����O��Hlc��2R~����^�z6I�C�V�ƻ_��&I�N����rP�j޴�iM���|�4��� ZM���3��vM8L�r�ó����˲jD��-��I5I-T�O�ݗ�jFO7k��T���)��K2ޱ�s�n3���ܬ͹T��X�c��yf����gJ6�a!�c����E��d���Ly�C�0�,�Qa/���Ȕs��4�ۘ�n�[��):p��8|g뿞٪\MI�@���`-�58�M}f?�R�_u	8x�� GkR�៮][wQ�����w6�C�2�(2;�?�W�����9�.�A��G�G�,L���S
ɻ�7�ݫ;y՝�	�"�?�z��q,J`�;m�jM�%Va�c)�����$}�
�_���hI����v°��@/=/�L�KO�7�\�r�7 {��o~hw��'.Um��D�"������?�U�%�+���5�9Air#a]v�m'Y�0�2򶆕0��"���Z�w��{V�3�}���!��<D�#(���r̄o����A�= ��e���.rrV�{�G������&��IZE�K�x��}#RD	m㶽�u�jVjs�+x�ZzGG1����s��:�D�{�']���`�AH��k���{�������M���y�'e}�Ze����@�,dT���e`i��y7֬�*ڐ���Nh�IX~(�N�vE���$���D�� ��Rò,g����D�|��A�1LI���H��@�ہ�X��핖�G�	ٮ;Ϫ�j<O����H���.Lc��DSҲ�E�W��^�'Rւ^ �5[#>	/e��L �#»������s��L����(%j�J��