XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��j�:>���U�w��Q�v�'o�sI6�w�MC� �m-Z����]��-*����g"-j��o��+y��zJ=0��#Z�0�ɺkC�p��D���؅�2��gxp�:� �?���<��\
��V.�n���e�O"�l��RCfP��ɑ�������E�f݂чl�o/���>��NG�E����$4s�%��A�nV��s���V���&�B��f�앜�q%sLz$��;� [���WЙn�ބ:�tKr8�d��
و)8K@5�\�?V�C��VME������#d�� �Y7�+��W+6�aF�JLĸ"s]r�5� l}!��5�@6�Yv/�>D���¸5[� �]�/��J%�l�Drԛ�`�O�p[�Z�ӽw�W� �;s�a.�G$"�5�5�\�7��16A��96��򹩝^�M]� ��VdS�ĥ���-����E�2���^ɬ��Ս�/�(f�p�) ��\����;�0b�,�D�n�(LE3�������S`2��EB�����_�lF|�?7��G|0��M�=4�@E�l������3��2d��Ն��Z�ԪCy��dY�"�د1�'�3�r˰�J@j9�Ѥ��dд0
����+�����o���
/����Z�b�3+xm��H�Dp�wB�j��%TU�A�ۙY�C)'"�\����'*R[W%��Q�J�D�`�p��`]}�GbAq�������7�R�h��n+� ފ{B?�ˡ\��o�r������Trٵ���5�XlxVHYEB     b88     3c0����)I�L����!+)�Ȅ���!z�Ԕ��ڭ_��[�B�������*�+R���(!y??��]`��5��Ц�`�/��S>�'���8V<��Ҹ��w�lm�4z��Ϲ"H�w&\� ��jWQhx��DnS�����4
T��\L�(���
��(��B?��C2g�:���.�6��:�-6G楻>i�~
o���rWq?�ח}��\{����U݊�1���ƾ7}BN�9/x�G�zD�\d�h��X;���a�|0�h����T�Œ2�����OY�_B�ع���u"�c���(��ћ@ �%\�cːF�`o��N+�ŷE�S��#��ahe���4f�Z�:��|I�&��^�>A�Pr��A�,U{M��[�/�Z(�K5��� �Ktc��,����?%��iWC~T�q�v��؝����9(mt���B�-�6���b� ��Ȇ�K�X�	�{*�Jݷ�
T9���0L�(G}һۉor�89���a��L�+c"���o|*n�W����*�6��~t��&�|��E�ٌ��� �	}_���'l�C��U��}���=��+�jy�����,n=�%F9���C������kml6:А�����=�f[7Q��g�Ѽ�^Nt�p�ow%�s&HkI̬�kq�^�܀;S�~�/�&#uj�"X�5�ыb���UVͳ߿#��X��t���s{�=mvkQ�d�����ƪ�{5�3�H��v�P�q�)�������4�'T%��E�~��X���ߜ�����p'Y-֍롫���^L(���#�łc2��o&���)�i��:�3�>"�T1��g��g��0�xٿw�+���3:$�V���]��e���2�G�8P��8��}UKC�i��}7GZ�y�h�J����� �X���-����;�J���͟>ww
�0Y70��q��L�M�