XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���:J�H~�\y⺨r���x�-Z�H��Q͉�}��/�.�>�lh5�sp��(3�|x%@����yof�vV�K�-�/U�9�1-�u �Jy���^�̿s ?���.=�~u?�M5?O�`�_uB���h ��yN�t����!m�q��FUNG9��A�ֻ��z��,T'��>�Qfð8u�
4��Z���ф��Hc��LnY�/k��a�\�ށ�9f���`�zH�q��C6�l�J}��r���m�dȾ�i��渒��<��bA���Ѷ�Oܠ�W�P�>�!}�ʱ����Ʃ��ϡЮ��T��8�wa�m2[1�(n��YuYmC@��(��h�	$�{���ƅ_������h���䰂u�R��<*�+?{#��RT� �MJ=�sMc� ���V1��q�E)��du�W�~ʎ(&C����2灊uu[�8̱��Ko��|��� l1?4� �ؿa}�s
��M�3���D�����	ϻ�4��h��k��~�h�~\�����X��UA6C��ݰ��
�Ÿ��0��ؚ�gRL:�����Pf��M�ڮmцf�*rRt#�6h��U'ZG�Z>��p��*�����@0��y�zD���� (c>HD� @�=�k���ܨ�iZ�Yq�� &�ѽ����6:h]�4�2��XgD!��G�e�G�,�S��!�o"|��P�D픦�p��7E����-��M9:�?(���M�mz�����vC���y%��5 m�B�rf�#�QN�L�XlxVHYEB    1491     490�Ő���m���-ǭ"���]k�Iњc���&)v`�5��O�����tM�0�O��%"b��-� �0�]�ST��Zİ~��}�0��3b��yxH(er�[-�5�2J��+���duQ;3�RwA��x��녂�^}��X��$�}JŅg�_�vP�C�#.��K$�:=���jJ�5��NHH1-Gő*n�:|8�Ym,��\E�UH��0���x�O��(0b�Z�^�&�4Q��R�]�KH�1��u�gu��w<CDAD��f���_�bJ1�[�ב�M?ėD�뇌�	:��Nn�o�o��+���r�p�)4�4�xx"�m<�X����oO�7ģ	[ZT/��w;U湌j	�b�o}Q�����'N2�mJ�����3����W?̉�Q�>>3��3f�-�X/�gc��/}2�[��vm� �%|�K��(��Ò�<��?~������p�@ �:tr_����S�Q�)��5]��y�y�l��qI1��d�|`9?G
���czL5;8E�:��Ο8���)qR�W��O��/ �J�ҟ|&Y��@'U����k�h$�>!�xM�j���
V�=�Q�G��Rp~h�"8�>1%
�A�}�4��q0�yx �v5�|����2т�`�� ��6F�0H欉���0��Y�qXص��E;b�ɱtA��!�:�~O~n�h�~r ���+9�v�����^m����0J[���a�`����q��Ant��m�-��hb}���GR�w
gH�d�������#ӕy>R�:
s{MGq�Ag����0�m�qn�T�t5�����/[�����a���j'��`HJ�l���}��\��m��|"w�Ok��F���0�z����|vd�L��1p�@���P��!�(R}��ެ4{�cX[��J.�P:1�%O�W��=��p��5v�Ğ�b��1����7���rBmڕtUj���L�ķ���Va��Y�q��-�JsN(6u1�<h8%�$�#>n̑�����yҪx��1�O�J)�ϤlJ��,L�zt���ڂZqτ�����8����G~-O"�͠�o��aA��t��Rɱ��yK�ࣘ����mPb�� j ���!��e�3���(<�1`	^n=���Z�;���(��g���