XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��FK����Qr�dd6i[�e(m*,�l	�p�|�;����aT+�f�vlNFպ�G�̲�y�㫠�)���}#s�g�P&2��դm���9�*���N�N��7ܐ�ߟljPJ_Ǯr2l��G8�֖K�� q� Y�AT6����$�e�_��"�цC�;�BK��S�9���d./�#�pKc�v�/W��Х���!ѐb �r����L^�x���.�� ��g�9E�J+r�m���5���8^d�s���3ާ���⚷�y�ϸpA��cO�K����~1��NΞ&�;�5�-O�Γ/A��
 �+��E��o&��C�xuS���t��6GA(����q�X�{�fl|���Q�z�AmfY�	2ϧD������"�ZҶD��Zj|�]9u�u���R�1ȹ_*�čk84h���"���3��ٝPޝ+D���}�r�JP>@�C2��+�Z��i��f[��)-�{H�ͧ�n�2P��0�5
U��N=���!��/y��~���g�Z�4I�k�(w̷8�E,�b��
IpJc[W�f��F)�{�*�����V�Z��R�M�Ԑ�����oW��ri�.�*���!}��� ��ZD�Y!�7"
��iP�U���Gi������ۅ2�(ok,�^�U�pUg�^�����	i��'���<���u�Q՝��]�_���-O З�]v#R,%���Z��d�Ӄ�f=�-nY��F���D��g�.���E�>�J��������XpZT7��XlxVHYEB    2fb6     690��O���wU*�@IT}Y}�����å��/��F�@��IV$��
f��B�\�2řS�~����B�eլ������M��[� ���Y� ���s'$�8,��[\�_NAC��©�5V����T͇-�
Z`��/H9]�l��7����RG��!z�H_�Ӕ5v�5e�)(�LN�����%YX|���]1$�S�_���� �Yt	m����jO�{���NF �$�Ch��b�ΦǍ�}Uh��BG_��ǳ���\�j>s� �Lw��#����h��q�S���8x�̹���W��v׬bh����6 /j=r����F�u\⊵#��Ⱥ�E�ah\��φ,:i���S��%�l��h��=�#[Լ]�=�|3#^��E�`��d��^`�oA�o,��4���O��t[PI}��;��=���؆)�Vs&f�x���l	�>SND��jV���eXs�=��@�=]��%�d}��%"�l^����`'��F�Q��N��F��(МE�y��qB�$y���k
)4���Ch�����,+P@#�R�����mġb�B�h�ϥd�ׇ�O�u��Z�Q�@��jF�O7�BA+���II�:��xӟ�4� ���"��������7��?�
?�,����� �\�ܝ%���(��;��E��ka�����B�s�}e��^s#ن�J���P>�aזk�~�o��8/ak6$1�Wq�i�1�`�� ƹ+�qC��jU����!�L/3���x�'���	zsU���~�H$|������d����W�Y@˄�Rl�o����v���#�H�4!�����BX��Ի��o�.�Ξ�W�j��8���B�� +\%{�kH���L.��Csb8��7��`Avn]ă�f��$�]�#�S)8�}�ΥZH� �
<
vb��� ]G3��5C�&u5���?S�l*�����H^���$J���Բ���_�q <J;IȰ�"����n)���,n�2�,/�S�$�]�&h��?ê��@��G���E�-B.1ц������xU�Jb]&�p^#pQ�W� 1 O�mP��������3�h.�7D���PwZ(������'�N�jA&i��9�/������S1j�+���]�Nݠ"b ��g}�hᯢ���3�&k+�Y)�N_�n������=��>M_�8�<V��yhX
k~TNs���0~i9��\��o�3�/����l]�Ei�.e��r]U�����$i��t�zt�.�����k:L)�"F:�%r�v��D����	���ø�c0O�%ّq:{䠘&W���/ud�0)+%���.�����n/�9^�m���-Gs���И�̚9�G�Ì����@��Wa��;�Sp���D̖)���o�5�fG�H7�de�Tg��.w�,�t�b��ܳ��2�ѕ��)��$�i54�W�W���;�֭��`�� �)Gcu����Z���6��~�k�y��wu���7ef����qO!(�$g���|�1��
0�~�� �޿I
���L�"1Θ	���I!_9�x�5���m}��vY�s�]�2���ފ��|nou=|����J�gTSb�hZ?o*�$�U�����`DZ�ͪ�~r��X�fS����o��F'�v�f�e�.Q�E.���cH�o�ByS�