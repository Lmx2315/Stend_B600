XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��,q��j9X�T���@����'��}�rp�q��T��i�h���z��m}f�nC
>[��r��2����Ȃ�kvO7S��C���:�VL�K)��m1���d�:�o�M8�t}&Β�G���г�sR���d-�4(��:)<�_(�*�Ҫ��?j����3�񐏫5�� �{u�������t�d�s�c�;�J'�eX��f'�_sP�����%�$��[]�*=m;;ĉ�Ш�喢,���(�P1S6ȋ��!���6��f:��̩��9M�*Ӱm�[B�榼r#i��n,�K�
�g-�������bJ\��F��|�6MYX����/b�:� E�˙Y�?��?a%*9a���������F@�c�VD	<�I�x�ۀ�݉�yc�~?�-��Y����ۖ�K����|ئ;��h�Ba�pY'Z�[��Ha2�S�I ��>%G��)D�m��slh6�Q�\X�Q���4K�<�<t��5�_��r� ��&WoZ?��H><��s,�p߱6���C|��.2����z��(��g������m�4�9�K�������Y4+���R�t���%"�Ҽ#���J\�l���q�N�>r��R)��}�/]�xڽp7)GB(�z;9���c`k.��_��.�~	LM�	�����ʀ/���hK�ύ��Z���VfT"�� �F�̋�﬎����@��O�s�mA��)od#�Ț����j<B��=E�1� %�!�FAr������S?��U�M�XlxVHYEB    5ff4    1040�r�!����8���U� �8�S��+Ы%���0���M��#!|�����Wl.�d�~�W���ߐ��o�v���t>�jӗ�qJ��G�<�w�mH��&�{����A-�h�3���#=n<�����h;o�ς�}?����κ)O;Y�	r�9#N�V�c8�}>D�IA�h?�~ߨ(��6C��	�ZTq�h��[���x01�� �M�!�:[݂6����F�5�BgҦ ��X�f�n���"���lY��]�)�	F���Ӥ`̨ʱ��$�����s�y(�!����jX�c�y��"�̱W� !"��C4(x}�K�(Q�Q~��qT9���B��=<�}��`o�M���0D�	��ꋽ�a0��=��Gb�=r��_��0���!�f�8�Bڙ��.Ў��������`h�^�9���EQ��8�w���o+���N��R�2�S��y�uݻ�nڐ��f�Ļ52�'eķ��Zף��H	�hDu��Jlz��vN[��:�f�k�2aښ�^��cc�<R��W����g��C�?	 {dw.D��U�Y��J1j�����0K�`gw1&��¥z���
�����]�sD�n_%#�E�E��8��ܾ`O�];�����Ttk�q���Z .B5~Oq�㪡�X�.����ztJ��INn9]�Y̎�\~n919�T����������ҳ�G�w�X�R�������r3�ʆ���pޝT�x�����j�����J{���Qc��2����,���aj}6�&�t?�1�0�|�rU��v=?���r���1�=�5���zHXO�Ô��6B�����}�0�`�&�8�F��l�������pw�����=�@�zIO��쿗�����^� &�%,�\PE������˴x��Y��TS����x�����H��40_�2*- �<`)�&�[)��8�l���p�Iǚ�_��
�$5�Djp��	��d �*��
$Sgh�j,����^�����P�S�+}i�j��r�������9ʖn/�9t`������6���[�c�5��:��kko��T�!�_o�t�4C{���<��ˤ7���cn��^=�F�Ea�(L��'�rS��bͮ��;��!��%n�P6{��W��өQ�Ycϔ�Զ[C���}0�%�ɎA8qL�k��<��N°�f����k8�TR�ŅƝ}���'����W&�Β��	8[�
(��H�Q/�p��j��Ƃ��W� دg	�zk��Fי[�@8 ՝^�*�����.��#'��iEv�\�֗�!T�C�Kw�3�,����~��b:H��s;�\=���cø�H��!f|�7�@3���q�"��J�*��^�h��~�l��'�+��Aʦ�:eN`�J�ֺ�8�6`�ߠdm�X�x�Hj�A4g�i֑���*�;3ӾHI��Q�3�,Dq���砊@���2��n�0t�q����6&W�2_ϗLRX��>��I���.dpf���4��M$&0� �:D	9�F���$3ӳ��[`����;3-7@|��xD������x�X4���Y������Pzȧ�@ױ��~�z޼���2}�����^��\A�5E��c�3wjA�P��m�Xb3r~1wVdT�� ����x� {��*h��buH���'3�x��>q?z��ɴ<��g{Ͽl���P���h����3f����ĊB/�����)�}i�:�bn��� 0��̜A[1���	���2�'�v"n�����~7i�����d���[�ո�&��.S��X���TO�4��@��!3J���ffQJ s�k{�I�:'�7w�sC��$|�v����!*�@rp �'��Vzu0���vXJk�bx��RV���h��*�|W����n�|���"aV5w8&"��v���l��R��Vv��uب��
z�y�R�T��[�76Q�H�僧��:Y��/h���|��J�1��nC�A���{��(Mz��+*_�Q![�_�����*xo��4�c��	�y_�۠k{�H<i �{�������T��f��a!��S�4��)�&i�ϟާ��sIm�"n�P�hHW����8)W�'���G��F3/�>*"���b,���e�Wu���\��b��ǔ��C����1�1�jx�^1����I�Y�n��W�@���8!WF�|<��f����p�	'Ʒq�������3��������!��@WOfΏ-T��:��ӍC_\�����]��$�/�M������@ww�xd@���h��ұ�e�}z,�Y��K5���@���;03l����)u��VA�n��<Xo�=U��ܾ+o/̜%o�)�x��I�8�6��i��+!��+􀀮~$�i\�#}xի7%�'���6�;�� ��6�Y"��*@ �3�����BԁT�n��G�K�ߣ��GgٺzXϠ�6;�B�n�}�"-Hvd&@։f��Ӌ������,.�1����z�k�s}�q�s�fA�ڃ�2�4m��y�4>ِ�i�Q�!���W4��+�y��qq;m@�r����u�	�Iy�aF�(��><-Z�(��r�'oUo��Je�K�ۑL2*o�]C;��V���Z^ԗ1�A��s������[�J�hU��P&#�`�⦺�������N\J�F�]<�k�����U�H��[��5/���E�3m������3��6Ǫ4����H�k�x�q)#�G��c�,5�ʂX�rOw�Z����X�=pS��\G�ރFy��h�:]�?�Y���l�,/�h�_8�����D&�����dXꀱ>?'}J?��θB\�O��X�ɨN��7�$^�q��P7�={6��U�+A��w��o������[���-Xq�| ���F�Y˯;�&�x����A��1�������U˼��I7�}a�8��Z�ІF��?'�^0���X�V��Cܓ�4�N�߾�Q��3TK'L�
%j`W9��bƾ�z��2w��?��?0
q1�B�=e���$G
���		��Q���_�ȳ�w��~Y��������?'2�sfO��p�{�����h҉�TjL	���ʁ�[[B�B�� :x�����R^c"]\��W�󥿮H�������c%#s�ZA��PD
�2�����,����},֢�ρ��1��~�^�dlq!�峲�D�(��E3L&�^���fB��~�{���2�5��B��"nH0���Yo�
�EH�mu����(�C��`>���0�轨*���~��1�3�Mc^�68��>��[�����'��,f�;S�ccM6+�Bǀ�0B#Y�ZL	{Ou����4��%1/���
Zs��_s�N�ʹ�g��,|C�1c��jf;��}.:�^���u��]�p����
IW�3e���x�P����
���<d)�6�D�t�]�QVÏ�9K�v��
X��N�'����a˭������P���H��G���M7$R���X ����>g���q����9V����Ω�!7�-okwCS%����moK��4r�6�Ƭ�D+�o:-h�Y�*:S�'���b"|_���Bd¶���Z��5�U���v�QM�?�S�I
�r7�>��U�FO�글���L�3̇쿥dF�o	��b/t�����u ������_W2Q�qς4��ǜm;���S� ��fGr}�T�S:-���彵~(��o.� �L��|��ou�4��*�/ض��%�޶*cN�ި"v(��i��QUs9�h��^��
�].Y���շҚbg�ٶ���ؓ����/L��!��(�`���{�����@�5�,�wr[9�ᬄ�]�{�zVeM����/��{�
ճ ��E�X����Q�ц�W��[���4�z׶�1��ϺH��j��6ؚJ��&��N�	b�U<��W�;fo�y|̽��2�i��H��W�I�����< �Uu�~����E,0;��[�Bu��,�]����PE�� �}r|N*��y���m!���%���0ݶ���إΨ�;nԎO���A�&���W���[ae���t3 �7��"����8h ��@p�>u����\�`����Y�t9B