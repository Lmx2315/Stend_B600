XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����t��]~١%�$/M+po��!�f��}�PEҿ�΋:Х\~�PS��T2��U�qԁ�ȩ�(���TR���զ!�^�7��.�)E�ٟc�iG�SA�-4�2���gW`ׄ�>�+E0ww�O *��@{rn�vX�x(�F`.~P@�%�8���n� W)���"�ġ>��^H�TpZ��K��2����%T��pa�wYs�-r�c���+�re�N(r>F9��r���p��>�T����!�o2b��gBA���zq�Owg���Y���^�=k]��( �r�8�EX�k���4;>���e"da"0<e�+l�$�٣��N�Y,�f��u�i���zr���xH$���z���n���Rw�9K��䎖��O�]3�g�J+Xqv{�M��kq0�쑭�T��c�'
����)dC��ݜ)�U��:x3�����:S�
9�&Z;��� ��7�\��%<�R�_K��z�}�#��.��RV����M��m{�?�Fti��27�LqU/��`���L�|4�:���m܁�*�7�s�Y�����_����{���$-�SaR�2���(W�/�(�>�%��b�kfh�j
�{f������b��Z�El���)�͇&KT�ƿ*$\�󰫂0�s#}A��k���C2�=]� 0q������v63��{�U�+��Z{C%:���X����/�%!m�Գ�B������%���[nu��}�,������ԛA�qXlxVHYEB    3c92     900��P�ҥ\]���L�<��7�gx�Ur��\��Jg��?���(��$�꿥���hz�&��#�����|�@T�+oal�ӿ���uyU��;>�c�>CAYyU���A덐���-���e}�C�=��]ssuT����[��g'5��w�Y#��$��@��F1c[�`a�/@p#pgq��n�[�������9M������A<��t��7 ��	���2'�t�<�۞>p���(b�V�	#-%K�T�����!�R�ێ��z�s�Jǒl6T�̻/��{�d��2�8��T� չb��Z?���.���0I�}n���l)2co�'H��� ���p��X'3[q�|�H�<ʤ}+x�K�X�<L���n*�5,q���S�W�����p�á����oU��c�Ŵ�,V� ���x~��[{�X�;�P�3s^��iȏ�ۍ���yN�8$N��=�W�"=o�h/�rP��E".��ãKc�$(r�b�!�Wu�� Z�y&��������h��.�:J4�r�Z$|f��K�׶�?P����:�I�^�<vf���L����I[{̤�,_�0��/m�	��Ɛ��{�1�zꧮp�_�r�*ߒ���BWmuʭi�[{45Y�6����e�t,�܌�6T��_�<��H\]D��P����B�>J��2Y�k^�o��%���ı�P��J�]|65�i�e��<q@b)z�:�+B����th`����`
H���M*��g�Y���Qe�)y`����32'��v��w����rۋ</�/��.A
����A�tO_c7�C�*g}�WЕ(m۷]��c�RY�رˍ_��������\�&��a�u���������������?�h򽬂ueە�XI_H�҅���5�K*>Ȝ� ��k�蘱�m�L�*#�ѵ�MVF"6�<SrM�y��pe7��h!R��7��O':Aש�YQ�@�ղ��+��/j�tP��e/r��rXMk���5�~/�f�+��d����;�|Xݎ��h�y߻Ȗ;'z���Lp�\��x�u��ة��SU|ˢ�# ���1����G^Pr�U�D�g"�}�{���1r5�#bK���́�r�_sK�F�[{��"�'����1m+�龜��Tߩg����e�G� 8��!��s���v�EM\P*�o�x�Sݝ�������:����<��>'��3(�k�$�5Pr�s��!K=�����U�A����M�%~���p�Ǿ���}T#A`��t&��/�[{����`I��	����2`�4Gb��n�\�h��jq�>��m�����H��9er[O��li7���#�ui6�� �W�Y݊�F���z`��tV۵�j�d�f�I|��B������э�6��#wU=�S��{,�1��~{����-K6���w�n�c�<�$ō�N5o�v��rLk+)
�b=��DV����ua���ٖ*��(EJ��):��9�(�l���z. ��Hf ��G$̈3vg�G/u����)순�_�=��Н
d8�0r�C���ZV�%�,�n�ٺj�^JUO��Vk�]uR�.�=����"�[>VK�e�NOYhe�
�4�߂����Z3�͊���{� ���'�~c%����S=T����Ё�,���}���r:�'D����R��SR0�+�Z��`�<��^�%��/���A�"���itu"D�&��qL&���� ;[(��AQ@MV�2��ħ�̴��/L�~�~�*���<���spME��L� ��:ߔ@�H����h%�q���j��=����8JEC˔��h�{��ڶ&�ʾw���.([_�86�ɣ_J���ަgl�F����G0�p��>9k��OM��g����o��D�G�t� ./V�+�k�`�����TFts�u��)��G2�;���w�h��}O���ݍd�?�Bt�[ϸ��3�="š�5[�*���Ӄ�E��tz�|������^�|�6?���<�!u:�#"a>��$)@|P�'|�>곱Q�j��3��O�\�}���6ƣ.����juV0t�0 ��$Ω܎���w���_�i��" ,݅�}��1@�b�� �LA���D���_͜t5D��+�g+ف2��H0�5�2y˥�svS<zt�Y�\#6Y��'�!�+Ș�}*���)�0�Q�o�X-y�����c�6��M|��bm��G�O��c�I.���AO�&�