XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������*'�ŋ�׫���L��-yG��S�g�;�kx P�q�Y�����dt��B�c�qz��B�>����&}�I�Óc��.Md�R�=���Mؘ�9�Ie̤���*��~�+���Q疻~�^)E�]��p��䃇�ǭ-�Z�F��aP��.����4�ك�ةX1z��??�O���J��X�'?�҇�E%���:mM�:sZ�đ�	C�OR�C�H�Hrrf�#ɏ��Q�a3���HKb���wM���]�z{әx-���E)��{s�ܯ M�I,T�/$ڊ�b����z���ՎAsΘ*G����rI�?6��u�ǌ��C'1�f/r,,�.%M��%�oEKu<#�ۥ6A�e<BsX_���J^M8�6�aB׋�����R��n�`�H!�wVt�=D�P�y�\��p��uq`,@ō"� �t1�'�5K<pH��9�Q��W_�b���`gy|���@��l�K����'OR7'��M�^�Sء; ���1�m���2F���!��˪'j3��b�t�56	��·��k�o���ln�]\G[��CF=�q/��"?*��G����ϓ=����pl�aW�S�J�l	❮�֤u6��x�TT:�ݼ�� y�?�x��ؙ���P@�o���1�#sռO�FT"�`Ӿ���.5G-�B(B)=[�M���_F�@铢���_�v
ǖ�^�4��媿�ڢ?�x)��w�B����rƊ�ۇ�k{.� ����*��l,���XlxVHYEB    7783     c00J�z�6�TT��rW/Y�3k��b�o�!�'U��8�[[%�R5$����	�����	�s���yC,s]B���+��v:/ie%�ڇ�Mo�m�(8=p�{�P �zs7D�̒ܢ�43�:N��%���*�՞qX��r�
��n��=(G-�i��I�}��vs_�
�}u��J�o���~��0f�1sVI�u�F��eF�*� ��TH�JP���܍)u�7�a��_+I�����8	���m�ܺ��JIbc٣���}s�v�Id�����_�63> �
�͉[y��u�K�e�$D�<�
�1�s�Ԙ(�-��C�x�g���)Ct^��*OxY���������g���+S�bT�$�%� ��`r���Bģ��ۜ�c1��F
�Gɩ��
 ����˒Xa��I>h;�f,�yt�+<��4kfƷ=�:'�ҿ�)�(@��Chu<
���p�B���>[�i�H��������?�DQY}*�K}6�4�
��:�{��FѺs$Ɔ?r��DXZ�,;��]c��>�D�FP�K�U�b}�}�P���L?�9�+�lt�Lb�P>������L�D��{1�#R:yО@�"�NG5��#��<	p��e��ӠQ@8;q���(�Cާ��I)b�Z@q���qY���Bod�����W���R"$C�\�[��$ټ3{`�,�ﳺ�l.lzs�7�Dx^I=}k�f�Ϋ;�v��lyLN�EɩY&�F�^��+`��a>�#��ZY\�a:�$�X�C�V	��;QP�(刚�˸MaV�Gy�^R������g*���>�֜N��فw���O5j�q�T��Y���L"Pp�p�w��w �EI1�ݟ�+ޫ[�E����9ae�#��B���	�����`�,}Д�[���P��;m%�K�r�����!���vO{ۺ6!�H���~���1����x���$I�L�f����T�Či�	I��_&����/˕�����U2���a�g���G@\�H�ql������@]�*ï����Y�.������hL���-FkƏE�&9�� {v��g�=�(cӌ�>?��1��1�z�+��&�SU*F�w��cz0���Uj�����"�i;�P���H]��{KMvp1-��)�nv�3J�p2แ�OE���`���w|�z Jb��z��#Yq��n �6�Xl(��B���y:�Z�pVx*�N��+/�.QH��Wm�P�&�݇3���;�ψ/l=A�(o��rD>P�à�bQ/�H����a�vj��cH�c��m�cVv��3�>N�U��&�F=���Bو��n�T��r{�M����7B��*��?q� 3�v�О%vٿ3@P��щ�%2��c��VU���J� u('j��P[T㩅�~~r��~��De!f�*��b������Z�3{�'��LѨ��p9�Eo�-s�j]�K��5&r/H���Q��>�y����I�����Ι:�ʽ>Pp�vO��  �B�<
9�F�D0/t�r�?���:��8G<m�&���w��L�V��O3�?O���� ̽���$np�~1�P�xT՝����,^^�W�����#eѨ���{l^��ރ*<痍z`K=h�������U���.|h~O�>p��+�Y�1�. ���a?���������1����!���96C��B���������p��^)TG�2�!'�(i��
-�wjE.��3��3�&tS��D9>�ӂ9��<!�5�O��冖�?Us�(�]��B��N�����S��ы}�/Wx߃;�$�d�%�	��>�عr;fT���ڙ_���[Z5����Ue#�SO��^pCZ��&�Q�#�x!#���E��4
�lW�Z��͈�J����o�	vܒ�+�
U�3.}	�`��	�<��p��N�>���~���ȡ�k��Xo��`i��m����7���S,�H¢�@Ɂ¥��e(	����_�"��O��ˑp9�S�j�/B�Lj����
%wO]�^vm	Zar8J+�mʜ�C�i�:ͨ07���˧��C�v����KH�묣����N�$��;��+a������|�I4MX���f����P�'�1
��z!H�qz;�P�iw@N������;��@��-ҩs9_C(Y��>��������m_��R	Y��F��V�p�Yg�pA��H~�#��L�@�`y/�G.I{!9��TX;�%++�E������׏��~���&�@��\���1	c��6�3�8����9՞m��R,/b���	�����Є����Ѩ�{��O��Q��O?=���<�fP)�"0�O�V���vygĝj�����y=���K.�2B�`���C܎V��1��|�ؖ&7�wf�E�'	?b	�)���C;4���������r�H%dy���G׺�W��m���	���_ҁ=u!�U���|iEmG-�O�n��@a��4}����s�ؽ@�SM�� W�P��e@��b�E�7����S��o��<���2b�mMI�����I�s���4��5dʡ��T�_�.G�R����sU�������AYg� Z��3f�Km�t�me�y�>��N²rѥK�9>MV�NW�ľ�E:���Z�d�[���1�8.��D*(��r�f`/As�1?:UB(��o�j[�ePK&?f���@ZZ8�5L�{����� -�.
;���0�Ca�������T ��d���`�$��;�&��@���]���9��S���K����n#����b;�P��=6"��Q�����#	�$��'�e�S�N��O�0p@6�RQԲ	d���N|��Z��*�7]��;�y��S,zP#�Q������^�ZV9���M 8��N<�\�}v:��QK��M�8����;�ձF8�i43��$Ǽq�M_�.ctn~���y�M���`>�a�/^��	Y�L��$S����`�w�s�;�I���|�8w�3�_��r#�E���y��x\C�8�)1$�