XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����O��S�� A�7y0��){�s��t��b8�)�z"�m�����k���1*���`P�l�5`>]�5r��[���ia�(���MGz�D���I�K|=�&&E��К�8r�vLq�� ���x'T�B��9@n��ؠ����"������Z��ftŊ�u��I�J0�D��gAf��4�JP"���~�ԅo��O�V���E&��8�(^�̊�#氿κf�	�p)M�(R%l4��	��}�U����aŸ�?Muu�3N��rp�e�n@�d�"���\4��z���W��ĮұҐ��´���C*J_)g�wֱB�j?ׅ��g/C�xU��<P�����)k�����Yb��`�2JqvS��<@����L�@8�_���G��û���+������R��h�.���ZI����L4l�M��r��^�R�PLݱ�;c��g��Gl�f��@w�n�FS��J��/Ъ�A��/����>f����*���'��h��8�{k��<9]`�����Q8A�8�:���{��j�u�x���l濾�>kuu�k�N�������00�Avd��p9Y3! �IV��:��A��f�UO4����y\sp)7x5����}���)L_ǀj&�Ur+ ��^��M�|4��6?C�>?}ȉ�v�6
3�k#ћ�p'&�4N�{/7�P9�D��6h}7�o�aI�9t�/K��x�������a�w�*a�S?�
��qq#w[h�0P�+�H��XlxVHYEB    1585     5b0]Lm�Ec�z�7&){<��s���e9:�9E.]Р\�ʰ��:<�6�`���L���p��{W.�G l׹�25��ygC��yP5o~`ڶ������B��B������B�m
�a��Z/��M�w㷳.L��N-�'��u�A/e�;ص��!*,a��u%QDW4�Ϲ]b����G|�X:Ǭ�"�[>'�~yOb���{�}�����\�P�$���f�e���G���m�����(�R+�b)J�\>S��3�/E�Zp�t5��{RR�!7��-�}��*޺*'���CKH�)�lv�lL�/�}gĩ{�6�4	��険Å��6c|ޟj���R%..�Q��V���y�	M�|}V�yW��e��Rd�j�O��!�(h�?�	oj��?�St��^�D&��b���E����z����[�w8$/�Y�M���Z@)H
�}���^EYOS�z�{��t�����D8g���t�A��$��}-/R���~�����]�Q���!X#0Y#��İ�Bk�7���g!r���>��i�Y�tl6���{�5y�E�ʜ/��j���Ր2.�E��<KS/�����l��Θ����ؐ"�v\ڶ����l�]����&�$E3�
;�r�6�� �RrW�g����$�	�_5���<&�3�n/�yFS]ˇ���`W�/�N����A��)�������6ao]�)��3��}�3L��ֳ���&�M.�#t��=e�����D䩭_�Եm+�����zm�Gg0�y5Ag�1��M��8E|�u�P�ɮY��4t!7ܭ�Ӆ����[�+���xV�����V9t��)���,���Ż�s�Ǩ~̳;�F��VKSRO5�:?�MK��L�	-��qm�s8A��@p2� ۷�ΐ5&��\���t���BC�F�n:5�oע�� y����w������S�t���w��g R��n'�G��*��J*!����>��­����k���>Z�j 7����0����$����i�M_�ux���M$�9��%��'I�fE4a���X�PD����N:\[���>��s�b���O����a+�<��\��[����9�/�9��E�W�i�d�S�W��a�٫ǅv���^��0�$�̈L����X�R[��Cau*�ٹ����S��!����zE2�F8�5#]���&\ʌz�6t6Z���J���UU�"6%��{NA�d^J$��5@9��������ɐa�Wg�P���O��8 �mhu �Y	�SF��2��F�0�,>�z��Z5�c
��W�P.��\4�z��pꖉ���ł�kz�u#��4��2�kUυ����#����ۘ�.I�(����0�N@>��� ��A[��@���4L�U��C2Cnc���e2��w�� �c_n�����W��9�G{Х_k��}�