XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���x�sb�M�Vh����7�dL�۔Y�؏��6��_�9�hˈ���;�Oo5Xu�qv���>L��2PA��Lp���c�/���0�o���,���� ����,�@��( <>�e��`x��k�}M�n�v����~FR�p�A񼓰!/�<� 8�9nڙU��Y/��_#�Z:�1�7�c	�qrK�~D.��C���6�O(���	b��'�y�LN@��d�g�s��5P�Qݮs�Ô��LB�{R'p]��q��|'�$?0��DWO���"ŀܗ�r硿U���u\�� ��>�����?%kq��$!�=wJ�9>+g<��&Q��L�z4K�U��*	��C #���ʀe�Y�A��#C�i�����p0�g��0W߮�1���Ok㤒T��'C�f��P�en��|"��E��'��^����B�,W��yyZ���3��+�G�b�nE�����E���
�\��u�Dr`m|iZұ��z�J��w	�v��C��Ӹ���~1w`e��(-����06����j��?,�ʈ������~^Z�W��2B�d&$�f�c�-,y(������V�`_U��<�1D��p�e��aF$�lw�SL�:>�HW�ЮS��9*D<��&=X��M���[9�FO`�F(��4 xab�.WJ�|䲱���K�F�0��_p���
�A�X0u�A��%�]��)zr�)Ӥ1?X��u��~�4�2��M��_~��n���XlxVHYEB     9e2     3307�����*�X�M�-̙B�k�<��0}�݂���T�[	e�|9�� Z/u��4�iVJ�U���m}n����N0?��k<j[��Vq��pf��J��ă$F_<�d�p�~7�_=F�R���{�a&���k�T��s��H?ں��̕����[{ܭ]<��s��^Q�X��6�V^�� ���u�s�f$j}lx�t�_+��Ph	�q֚��|eٌ�q�@P��0U@���2����_I{��\��6u�F^f�W���U�A���pR�"���y5T�rov=�G�T�j.��\ɀ�f�۝��_XKH��(w��;⟰� u��� J~�=�vE�)7|�(�	�/]�UE{$�f�p`疰��F~/T�l��5�b�Y��>roK�'�/󂙂wY���;�6��K~ޘ#���V!Qv[lFbA��;�'I�'ٴ�Z���["�¸6�v� ��S��dz�,	U��d'e��������@�U�>=�ٞQ&��F�#
�X���*�о���i���|*(!�H��:R�u�d�6��w
����ECYכ���5v'��i ��D]����3�g���~^\�D�7Y��z�4T{��n[u�v��5����p�z$���r�Zv?t�JPyQ���V����*Rł1��>@�!#�O@��*�"�~� @�k}|+o�����6b����"�M�����|f�9;�h&�R=4h9�:��&i�T���EIv��a�SaJ� ��i%�Ւ�L���=�*���\)�Q�D���0��*�퓔����e �t�&�b^<D2[Poh�������ǜ2�X&�9��0@��[��lj