XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��� C-�aI��B*�����^e:IT�&Q6�c�i��CK�L3�H�K�8���b>�B�&���(�m��~��3b�}��u�����hNW���.߈#vh␉����~�+ߝ�&��iO$J�D&[�D��{�D�N����W(�R��	�g1h|��JI\��c׼��"�`_ed46��X���m���W	xJ{�P`m�w���$�l�Ǜ�(͢^��ԟ,���ӟ��{���͓��^J�.�4 �0��M���������+��H� ��.9����DS����Ul���.�|V�=�N[D��gT���ˬ��B\���
���5\�Wv�,�I��h0� ���r)4RP�@�	\"&2��%2�wR���L�J�U����YJ��D��̀�u���RwzXǝ����p{�xø���85�����T?���� R�ll���F�8���5T�:ݑ`�q"��`�� �� �D���� ��<�I�]Jf^�ݱ��GV}��ΟF�Ǆ�}7���}�Ǘ�9l2;�6lt
����:1��y�k����0 M�"����Xn=�P�	d+�2 ���������ό�祧����n9S�� ����X�"�8u��1c�p�0
�M�%�
q��׸S%�?��Ơ��z^)���'[���&Q���?���ւ�p���P��H���d,f'�� �����2�읃��W��+���_�5꽍�K�y�wN�� Ca� �|)�e�x)�H=�v'�b���+���}��`]�2{���k\XlxVHYEB     bbb     480�*rO�	p��$��K��a4����3�~��銸�F��4sQ�6�n�/���0�Η
98���H�o�#j��df	�pƴu�*�)+�xY�w���]�L�%v.<�1㨦�[ǫrI�[��b�@�%�1�h��hG]r.R�Ώ��u^�j{}Ű6�b��
���v����J��E$+,:�T+��]"�0(\p��)���=�T���O�.��m��g���-/�X��01%��I����&&���;��с�D�pg�Ts0�t�`w���\�G�;K:d:��
��uկ@�
����4u��n��'�W� H�~���f��h�|c��q��y���[d�}|�8� ��Z=�篶�Z�6��ʘ��ŧ���3��~XM6/�1�D~�O�;9�h��b�8��ǎ>�D�)��ו����:utuz�%���7&�m��_��.�-�]�d4�MG�EV����K-If�[�d޼}^=���A�k*���<���5H-�_Q��(���^�,B��3��a~XW�� �<c�+vQ�?*����_�Y�N��b��Z��Z����/�U/]���x�I�P8nV�.f~8��7�ݦ6}�+���"r9�S��a6�H�^�7*kF���+1D�,��vo���q+�%)&�y�bx
ޒ���$?��s�����[_1�K�i�C3!�Iw�%�ڀ�{Zֿ~L]�~[�d���מ
��0��Q� �
�	�w�� ��ME�_G�g@)$��A�i�^x���)�UI�-gR���~Y#e����z%Y���99�d���	]���� �]�u�j�|�Lx0��8U��'� A�O��
���X�us~��~�daR��}��Si��?]�s�FDYT�ñ ��t�"����,XJ�0�V�,�4*�IJ�[��FO1��](? ��������(�y+��p�ѽ�I��Zܹ����S�5�������S��HJ�}�d�R�|�����i�3�i��V��M���-ֱ�`�c�Dxi�5�O+_���bHm���;�A�����F:��&������acr���/az�����V���(��@Wb��N[�n�f�P?���F�:F��cP�pߐl�p	|T���pG�>���|/DɎ8