XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��N��].�����A���O��$A�k���2T�_�4j��:��L@"���(Se��"9�d�BfcM���^Z�������iޛB��z�)(�:��-��J��I۔�]��Aҁw y���S�Ź�P���� ��_@n^fň��6��@��G��}n=/L� N�a[X:8��B#ׅ��&�;�iƜ�E���7�;O�����>[tA~�O-$���9dw��m���~V �w�wX�/@���Dcf������h��4t�^���lu��e#ϗ,k���mqK1�Ъ?�\������'Q����u�$��+���Y�uSQ�,.5-�(Q�ͭ�}��@�x��NL��������,x�ט�B�����A��T���bO�5;f�k?A�����4k[r��O�9X����=�P�a������w�I��{�/�k�W�䣠�����R��*�OU-�0��n<|���p���@�*�!�5���5�f`�k����b����t���ہ܃�~�ݑ=D��#\�KH����I(�g��J�2[�a+c�A�Yuk:k�sJ}y{U+g�b,�s���k	A��������/���闩Y�Pq,Z�r�G�Mz��w��/�Z*�XD�� NS�����7�B�"�rj�?)mD;]����QM����:���-�z��tmL|24��[n�CW�Z 巒����(�8��R�F�xs+�)py��/��S_F�`Z�TZB������F�@�ߠXlxVHYEB    50aa     790��c�UI^n����؏��0���7y�;�I����SkiY���r<����W���(�k^Eo?/p���	5$:p��q%�y���4�š)Y ��q�__E0u�ȆL�$�)�C^i</�VR��kx�y4��2�մL�����*Y�b����6W�&e8������\91�"�m���qr��L(�a������Kd���gO��2\���1?\�!]�e��Z_�.�
}�O$�V���O����y��Nu4�z@��W"8x-D" �;G�{9|���S�����̊m� ����bk��9���V�zZڗ>���g���ch��t�$X�p�-�w!=�c�h�o�=¬��$�|�W7�d݃�7:����_�uaƽU�I3����X�����x��"�H�-%�����������-���B�4�B�3M�V�'/=j8NBa�,�~Pi���C���f!lD�"0p�s��2"������)=�/zx�p&ie\20;/�s�
͜My���)a�~Z��G��vJ�gӥ��Ѭ��XQ��)��Ώ\D`)Q}�o�A��d�6�5*�ؐ�lE�$X��b��ݓN��Br���ivM�����Y�TMp�"�3Ǎsc=�v����6'�k�R��.f�1�]��6'u�>#;�,M�*���X��VHU����!�]j-=ҷ�iM�^6�Z#��S���c�QaY�R>��h����"|�ADJ��|����.Ab�\÷>�`�0;0B�7�}̂��N��K�6,.l�}�u�e!�t\��&��ǵn�)NDxBVArc߃��6�#��>V<oܞ@E��Tɚ�.����5�$R���7��FP%�I�B�4@&�A�D���=�����열lp�'��E,F��U�x�J���	����-�NI	?�qH�_NB���E��ݞ]o�a�X�}y���k E���3Ehښ�G�s��˫�D��G��]�����K������^�H��Ym�P�k8���x��:��� Uxt��RhtL��b���~P�;V��.��=��iB�n��O1�R�T@�/ɭ{�`�@����^y���Z=l�}��]���xX"��`��W���쥮�n:�RPE.�HN�~Ln2�K�򩧧2�:Ab �4�C�$d�o�E��2/�c�F���S��{��y�ӷ���y� ���+
$�u�ᯛ�rI�x��y�-.�?�օ��:��eR2a���jd�r�*`��D����г�#����w
U4�[��D/���9��{�%��"A�+��K6$O��IH�%*��m�z(�N����CT�R$����vrXlM��}ni�������&�l??aˉzS9z@ض�?K���Ls2�4�ƥ����yj���;�Vw1��b�7�2��}�2��l6�I�e��D��w���ۭ�	]�������ւugцMq<�RBjc����{�G��y��2��sL-����(E1A~��)ɪ7<�):5����Łu��*�;.c|Ș0���B;�� >w���u �b�	A�AGY������'��6��" �<2x�Ԫ���I���~�n@O���&k�3/����7�M]�C�t���N8X<�5�账PƵy�i�7ő��b��훁͟��h`� ��S���+�S�Ax�oI�i���2m(&{��� �n�<��=�e�U�M�HC=��z�-5ƛ.�`�1D�	���&�s;�UM�4�%ʱ�9�z�9٘[�}c�R�����<: z��CGt"rb丑VTI�����F63����A��ѱ��1K���	$:�<�o�ϲ�R�Fn��'�w�WZ��⑅kwè��x;X��f	]��� ��PR��8�4M[��EE-(-�è� �.}Tn4/�_=wܦ	�)e�ܪ׭�M
�����/Pǂ