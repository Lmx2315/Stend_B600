XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��y���W� *�A���.�7���誮�ڋ�+�r������^�l`�X�+�e	Ń�'�#;0��ͯ�v��;	[���K-���0�BH^����&�EM��|3	V��B�z\���lϬ�
l�.U�]L5��[���5ci!��ن3�߫�E�_�Eg%w��ڪ�<�h�g��(D����g� l}�c�'��3��.5<l�~VS���Fбu�C�	���<�}��{r�q�(h �٬�#a�3v܊�s��7[���b�Gp`���a�_e�兎d/�GhS����ݠf��a/�4)E��@h�tj�o�m��&B ��p�\0�s�� �=��hh�I�TxI�iSz���%Bqm~l-ۺ.Ȁd���!.@q��F!�2�����,�I|����]�a5ե'�>�Q�JH�J���� A`��G8L�-�:g;�4#m��l�:�,���N#�#^�:n��E���7j��u�E�KW"�A�e�tiy�6E>�ŕ� ��g�T�NP[��%]{�֎�9�G�=�2�����upw���a��Յ��Nr�"���W�0�����^H�'��u��WRW���6M�NG�y٠��mtt񒞻M}ׇ���2�跟@=� *��H���\!8����E�R4��g�(ۻp�-*���&����)�!��dWjѸz>oBM��>Y߉q��r�]�ľ��MS����34ꁡj�� 7��k��KT��9���3�P���V|�����V1��C,�J��m�wm�J[?����~b����XlxVHYEB    3a1c     d40臼�U����	ʭj_���=7G�T3�f���B	C��\C5Y�G�͝r�q:ȥ��!���C��@dz�Ān�?!9�V<W�IpVZ]�J�����]���R��UJ��8p�屮�u����j*�V�3V�ר�	"�.�=�l��d����}iw|�����������g��E���_w����޴������DD����y�/�X�;���><Y���
��P��TyR��9V.s��]:�>���_ͥ?9�kH�R���X����N�E�n���<tLq,H��G�!�Ze�e{�9Q�V�GԔ���3!#<.�Ptaz��2xb��;Ba{�=B�5��h�b��k ��v�ו��
��\�#d���Mc)�+D��>�Ƣ�K��P �8 �%�e�M�U�z=e�� �m��E������ځi�5����t���wi;�=Lp�`����ȳ��9�c���������9�"��I�P��,H@�9�[��F�� ��ڶ���\��}��/l�D�v�Y�;����e���.���W���jg�r⩓���c6f�@�Rs����0%|��w��Mm� ~%K�?_�Ȍq��W>�s�65Vn�:P2��l�Z��8Zk�#��9�S�z&aտ|���mx��z|j4���-p��ũ�*��2}L�9.,Z��`e<f�lg}��@��>�s Rg(���7��u�0 J��E�K��r�ڿy��:��J�_�M�]4`u��E�Q.���5��<+2f�I=�2p�)�v�Y!^F�������HV�[5	4������'r�{�ζ�7����_��eo<����?��.!���E��~�[M�1���K���J- 8f��7���߲����&�a�N��߀����R&�S��"�C�}}�U�'�e��LM�A�U��:\6.�ʝ�Le�*���{�]��B���}y!�9�t�/Z��A�b�0��V��MΩ|�,籺s�{���F�50���[��$�90�i�ٺ+�F}a�L��n��V�zzE��u��l��ו��,c�	R����y�v܅�����FHD�������$,�H*1��P*~Ì�LvU���N����t��'ԁ��jL���@pH� �.��.B_L-H����>��X؎�@�b� �: 9�����f�˔�S[�wgd��,��rz�.��}]�ˇ����c��z�`�ņ���g�,@h4�)\���\������&�-��N=���������l�B5���(�R�9�FCu�L���o��_�u�S)��T�V��`��p���k�?�:�p���WJ����}I �� ~�AfY幸��+�p���}6&��צi��d��Xq�.%QXI�Q�����G��c�?�4d��s+;�!�@�-qa��6���cy�X��g�ɢ&Oͽc��GK�(DC+$��������[�T �S�� �'��Y�A��,CiA��K�eQ��(\0r��������y���V<��y�^�7k����g����j	�Jl�\�1q����D��,�ڠ��Y�7e��_�0G`�Jog�5�q���277	�_�4�B��厜>l��n=O7X{E*�随F�pTe��b\;��s鮯>�EDjIv�9S	h_e**؋�3f�j{M����
��'ȸ����o�9�G�U�F�4.	�f��m/��ݲ��x�2Â��E��y :U����U�
o� ��VL�v*���*�~pͤ_����U�.��_�T2Su!4l<�=Է�?��Tz�R;��\�8����So��QD��qI��nc�(�c�'klEͱ�XR��s�sa$"7��?�N�B�M<�u�gǦ�{AC��V�W�gR-|UF.�z�v�8�%#d��D�֩l�`��f����3T������m�TXI`BsD���%ZVQ� �a�}W?�E�D�E� \�V&������&��a����cQ�=0��0'ȏ_���1��X6m�v�Z�m�Ts���ޢp��b@5�?��|��*/sۺ�D%$_\՜�m��E�n�����9�(�c�"�'T��g2�R:~IU���~���q���b�0'��X���@���႐tSW�����T*>5)�Kp����ge��(߆(L�O]o�֎�A��jO ���a9�0]+'Z֊ @Gf�p���GJE�M!I��F���FF���������ydv�:�qT�	"w,�䤴Ș�e[�咂T[��S��:b���E� `a��2�3�	Lur��`T�?��3	]�����Dy뱅1��6���MbaF�`ը���Zd?Ǘm�R�T�9��|?N\��:����Ώ{�l~1Q<)�&�7r?2.k�,�@Z��M
��)8d�#�7�c�^��R	_��L�M�����Y���]FS��Dn͝#���t��V��F�<�O;�LTC�f?�J��?*��Sy�4J�ɘ5�	��d�AdeX�o�[[��.3m�pa��o����Ӌ��،��g�|�pc(V&ti�h)z�S�Gf;�jʝ�Өs��$��X�z���nI��'�j�#�O��pK� �q}�F�2ܩ�+$����W6@N?n�@R�(�����x�B�[�\���Ɩ�,nd-��&?wߡ�`@�j������:q<��}�0�H�O���	�de]]�C����k��(�+��"��堬[�SY�ا�D#�E�����������i��(`�fL,h��3�^����@�!KR���qո�:s*�����W&�5������̦m�h�\>�h��ޘ�/�����X��G�Y��w��jr���N��H3!ߵ!�;�ek�Q�e'w�;��R���"9<��|ܐl�ؘ����� �]����E��aEd�d������,e��(��?��!=���u�6��Tϲ),������6��7����wc�7|`�9�����ab��D?y	+�#d�m���F����W����ϲ�h~��h��:�Y-�snn@d �U�j{�Br��ǫP��D�{��Z��@m4�����_��(�ѭ�;}�F?�=id ��)�Ҽ�������4;ވ�>F�A�ƛC}6�SA
 ��B5�����w`��՜<s����G��9u�]���.�_�籃)�{V-#l���v�Bay����r�ɼ�&^�-]՗�rL�O���\�tC�.�v��Ns��&o�#�ʓn��v�szځl"pG�ny9�FN��Y�vf?^F�(��>��  z
�±�G��iw���*�4+_q��s"c	0� �2c�{Di�f��1�1~z�QJ��x����C���I˕#��JV�A�b�Cm�Q��i�ZPr�P8e;