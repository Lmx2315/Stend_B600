XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��A���]Z���'=2��V��SM��i�jz��*�z$�5�]z��Ł&w^�����ċT�Ğ�������{j���
�2u���/�����/zw/�K��0S���yTKlNׁ�F�}�OĮ��!�MV�X�h&��X��R#ԯj��qxI��࠲��s�4RAG���=g�	�� ���	H�M���f0=��H[ܧ�"���m
��V ��	�����,�'�R��
�g�e19�Z���4vT��FQTкS!��D�)����>�[�:g�yH�~ȕ����,ʮ��{��ݶK������؀=Ⱥ��G��|?��UP��樟��B~9��I���:� ���Mz�2�I����񿗕=A���JCa���Os���b��4S(��PB<<��st� q[x^(�pռZ��7g��c�0�J�Պ�<9x��e�n��ј������zNưJ.�7}� ��i=�όJ�Pu��'5�Aq���~I+A^HB3�����z�g��5g�j�ְ]>���e�m�CH�G�*f���.�}���Ŝ��DQ�ժ���,H��D߬,�|��.�K[P�֡K��'i�/��hVJ����T���	д�C�������C�������)(��ʃ�);L��7승6��@�v�zEF�f�`�p���P孞-�bqA�(�<s�ߝ�<��k�ù�Ь����Hd����ÿ����'u,&��Se���/�o[n�~�%�cxk?@W������XlxVHYEB    7738     790��	Gb��Ш�e& *t8���3��6Z��{�U����3��Y�d9���;�5kR���o)���f����쎢%���jC(7�W�/�Ni�Å�O�"-t>���&Kr���}P�y�m'rL����]��9�+	�Z���;�m�EU��Xh�����Wr���o���X�[G��֓��U	�Y��i�Nd&�Zf��n�c�@��E��C�����C���c��c\G�H5��`+4<}��Ɯ�3)��Qi
�� 	;�l��
E�K�HWr����|��y;'�郜=�>��0�f>���h�֮p�.i��K�@e.ZB��-��JT���N=��Z��<�����\���S�*�=m��٘X���RMİJ�s���ǋ��#rl���x-�m>�l.��(�jK���1���eORM�U�	��*�����Mܹg�c�23'�m�7j���Q��9�:s�cK:�r��G��~+�M��j�0�#,�M�r��N���o��Q��z����b�2_,~��9O"��:��m��G����}]�4YM��+Zѐ,��!���*\�]YΛ}Y�7Y�s��m�q�w�9Bɧ�q�\�F����bO��"VY!�j� ��`���!,S�!ƥ	@�w��M0�p*�j�� � %�Y�ukݻ�r���-�f�8Y�|W�V?<l����Y�>Q�����y;���J����8�������N���b���HŜۦ���S��[i�!D;06W�m� )���#v�*��@HF���������r���}���].��S��,&�o���0��1>��58) �tn��6�l��J�jB£d�*��p蟐�u�zCT��4�;u�*u��z�6c�yAʟ(�孃�CҖ��^z�:@Ƅ�W��ש_���4�a�|cG�^b�A�p#Q>(������(/I�'����C�G.Cܢ�4������K��/h� ���!ޒ�z�`pj�N"e~��NL��v�vZ��Z3�]�vx�nb iRhT|\�!e!^���id��v�畈M�f�Z�(�- :1�6Ss��pH�	ޟX��m������|DxT�%�8��=5�CB�����rN/�c���U�@§�����Wc+�w�b8���/���}��'�<�|47@�ϭ4/U���ڜ�	��%e��hc�x}ӈ���Gq��9k_Qxo���fq�R�BqB��RQc�T��f���*����^{>Ė;���?��TT���-���mu���Wa��{T�Pe[I^�*�s�j����/��o[
O��+"΄-�u5�Uq�?6F�w��z�?�s��t�>mw2�	8�>�l���[� A�ӐLYu+���<:��Zg��eg���3 �e�!��aIB��*׏S[	��-�h���U&�WÖg���P=�\��>��H��$ó�}&8V@Ѫ�s�"�~ȫ�M�4Q�>Ƣ�/&�.����m���h�����hrs@,U���U��g�),@�TV
oX�Qa&��i�t�:���~�t֓ь�M�����8Xb��!Ws�*Xh Lp��+YǗQ�J�O�A�߲�������2�����ԙ���F�G��)7HY�|��$lj�+����L�Lcfʡ���� 13g*w��w����E_�H�t��f��m�~��\M0��t}*'��A��$#\v$0`@PG�}��|�E�-�q�$�sX���s��wjT���A�@(6��U1/A�)�0&;��Q^���t�����{�v��U���<�l+�v�e'��U�h?��N�֌tm�/�%�Gn���CD�V+���%l	({̱�O6��"��vtЉ�Y1� �Ȱ�@��U���P<�@���ǉ�Rz ��E z�:И�^�sD�.i2FV