XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������ǳP�a�h[�:��mx�q'"�-t%�Ν:�}I
�� O~1JD�)�Fr�s]6Ȫ�~�����?�J&�2eRHf��s&�Iݺ��Z�9tC-O�'D��>��_�e�N\�t��|��=�[��10��^����d߹�a�{��L�,�#x+����^�yE�l��(	����"@Ԓ/q��i��H�-/����k��
��L����Vum�5�:�louD'-�n(|����]g*5�-��,ɚdqu+76��g��c�-�m�w�x��xE�!�
����=`���G_�R�9묘*(U,��p�L���������
�Hy���$(j����lG,���@S��[��x��4� ��f���H�$e�h�u�',ހV`�kǤ ����^TZਫ਼;���&ꡤ��@ҭ!=�*x���h��,�|���Nj����n��l�c��	���3n4_A��Y���^i��� ��;���`�TKW�p#_z항�Z�Qt��R����"OH�}&J$�O�(�Mn�/`t�W^�57�3e �2,W�(ڝ�O�9��R�I���_���f>���L��H�S�buy�L7���͐p�wZ��e� 7F�����YU�W��nY�����'%��fڭ/��_�7R��b��\`��A�.�ύ�!�bȳ3ih�#�{��W�"/%B?��M��=�G��_��i�i!�֩xMwk(�����Nl#��_�/���L�x�kt4�JV����H��K�?ad_nXlxVHYEB    41be     c40���\�aٴ��W��Or���S"w[rd��фE"��;f���y>#""��_C�2z[���h�Ѽ���[h�cgu�:�!xg�:$�XSG��YX�#�(�W��ޢ���f;��i䁉�bD?��e�]�
��g���36�N��������Un�9�>l �ndf�V5D�_�ߴOLqn�X|����V�����f��B�Uz��7p���YM��"S�4�E��vh
~!	#���R��(v6hzf��|L_ F�ۃ:Ǖ���U䊠���O��W<B ]h�x&y�=�V��͗`kZQXz����;>A떻���R��v���<|O^�>���"�3����Fu'O_9-��q������N��5������+� ��_J���|I�KNs	��@�&nCކ{	�"����pВ��:
6h��ȡ���|iNh�Z5c�QA���7�;��xt�ٹ�9�\O��L�xOB8�rE����k]M�e�\��0r�؍l@���^^�Ĵ�����<���q<�����C0��	�ged����}�K�g0�dfd�A�վ�ȓ+�=�>e��Z�U��<C�ٖ}m�q;�.{j�Ҟ�͈���擑������j�Ҳ�ʍ��iP�9%v�?�i�C�T����^X��`�k��毘��ƍ��R�S����,�y�Zޟ��֤B�J�f��Иݪ�x���F���;o|��[J_<��|�4��Ǚ�iq,��'�4DJx�M@[�J*[PU�?���w��8,o?Xa?&����ԷZ�
�D���Th�,u�z�r�~�=!`��e�E6�X�\\���oqo�]��b=�O��썘�����&��"�11���cC���x�=&~�Z�g�ܽ�X�Q�;M��c<b���M�H��!�9ËO�����/c�.�@4�-���Ϋ>��l�_E@'9k��@:PP�K�R���V��lIܼ��Y���I�x��c%���3��c
iw�-�� R5�L�k�eF>%=�`��2�^ۛ��[��@�~�/�/`������uBr"��T��|�ȵ� �@�@��[�\ɌF��M��+B}��Y�A��0x`˸K�|�.��GsG������W3ؚPԕ��>�C� U� ş�%������Z$�&�Ed�
����X��A	��.;�c�!��{k˙�}�^-%�Zp�<�[U�[�IΊ(����%5I}��$+Պ�����>l��jq���-�t��?ʨ���}�p�� q�����Hkٺt���iǘ6|&ͬ
��G)�-�սr��ɗ�M���y8�.��i����p`�7���[�Wf���Fi���;&�H��9�]���@��S�o4�cN�f�e��+���lA�Pt���υ¶�bͩA�$	�e��.���f��|r�l�u�/vGS�Zl�zBg�'X䛍1�f��dK�Cx���{o�CT'����Ceܝ�U�N��g��CRJ[A��I)RQ
e��؞h��W�I?��L�f#�yL���$�x��v�,M_��\����y�i\Ha��Z�,�����>o�;��x@��
|����������*�`^?�pK�#�ۻ��
�9�Ge/M�"��ŗq3�MZu^a��ʇ�A/�s|�<��\n�Ž���l�7X�]���h�� [;�T���g��bJ�+Z��x���m*ơ��[��αkv��!��X�C!�>���r ����p9`W��&Szk^��QJы�b��Qn��f����:�b��%��Y��*�=�,˾�ii�@_���G�= ����onGl�X�?	��q	i�59%+�G�����]~�ƄkR�S0&�ǽ�<Yc��q^<x�˔�57����d>߸F�,�%�$`a�Yb-��x�V�Gb�b��l�Z9����D���m&?�~�	���@��&涴xL���_���l�܌�P=�[^:��ΆI�x��-�����icth��f��D�.�I�yG���y=��J�Pی�/xDq5����j��.��Q�	CO��K����` �)�bA���!a��qq���2^��6S;�3��*���\�����������BZ���U�S�j1�1'Lnel�`:x�T��{���"������
���]�/N�GJ�6Ү��~��D���=9�Ww"�$5��\�r,��3:�V��Z�/U��������
f��,��fvU�GE��<RP���?���Xe��������u縣�s�H��K.��eI�����p�r��p���ͭwn�ۓ�$|�o30�,��g!Z9!^�ʒ"�֖z�l���ƪ�]�^i�y��d��g\UH�,�r�Ti=�A��%Bz(�x���� I9��`��N���OZ��@�Gv0h����0	w���aٯp�n<_�¼�94��/�z�c��>j�5������������M3��GQ�0�\�W�O���U�;���&��cO�����6<����S#����f�@��MbDM=��<p���Yn�X�D��KtUW�%D�����'Gop[���K��lA~��M�>��ٹ�qb�-I7v �*5#c:��c���j���)�/�ԢpЗ꜈��Dt� pⱇ�`�'��'�e��Nu������ ����dD��<�_U�Fl6o����VG4�ԠȎ��d񣏠:B-t��j��Z��a�:�X���@�3��N��MR�l�R��%L֭�N)�Lt�8Xt(N!q:#�y¸U8��w�D�tiAW����/1;Tj��ﻕ�3v�2'k�wYZ���F�*|�(~��E}��Z>��amw]"���4�t�۸�H������KX_GD2���`�݈l�W�!k��q�x��Wr�z/a:a,���,��p�s�� V;
U��9A�����W�g�kC>c�X�Y�`�sU87.L����]2��6G�h�p�f�ݩ���ז��h������j0��<�k�4�B��l���\ �6�X&)43 =�;���l�
� ��+�+W�ki�eM��|�3�*YL���e�+��o[2��%����׾�+��{���3��Dk���]ÿXΘ"�#��ˬ�