XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��� ��b��?>f������7��}�@a�;�\E��|�z�T�D������)a��(<L��"�AF�����Ø�:�*!��J�^ \�چ>��4t�<������eĻ�����-	k�t���	2�?���8����Moq��B��κ�~��qBͦwTjx��Qw��{�ڗ�����ϭ������[�w!��5*�(H1��Ɵ�3ѝ��R	a��O?C~��MU>���&�(�ڝ�}Zo��p�%��Q���+���݃��b��h�/s�����h�3�j�!���g���{�Z������c����v������UYn���#D���A~]�=C)t��|�h�-iZ��a�P��On�Y�-Χ ����Ϟ�:�����L\F������3���aM���CJ_�b�xjJf��e������M��C��Z��]��_�>6�*�:�m��~wY8s����h(^k��^��5��xz�"1��iQ!,��G�u�]����*�FBw��uhMg������U���O�:�'b�����Iy{��_����!M�m;�{�D�1��)8���@��U�#����䦂�� Y��z��U?r5S�9�Gy%Ba*�q�JG���rr[0pg獃�F��9a�B&��C�편�>��ُ�~;[�T�F��P�Q�Ѥ܃OM>F�����+W�,��H���ܕO���tStZ��檀N�,��p�)�=�I�7�qWv�k�@·��RDJA���ɱ��oXlxVHYEB    6fd8     c30���-#��%j�I_�n)��L]�͸p����Uj[�.q8J�`	��w��>�xK��p���ƻ;Ȉ��7��<�	��("�z7�ׁ�kr�ܨ��'�u�O�(�W�z�Y?*F�$��+����t(A�Jj�d�6���U熝ܞ�z�0m(I�$C�����0Lq����W�l�F<I���p�ózmm$DH�{CS����]�Uq��1��G�'b�RF�)�}�ѼGp���~��R�vJ6��F�{�`�{ǚ�C��cT9��|�a��l�i�s���;�#0���#�a�Ah�`+ޭqH��\���5F2��,�Um9�̭��tR$g���.)KU#z�4*��`�Pن��֞v��޸��Ѭ|���U&�X
��Ф���&��B����f����
'^�to�������=���-y	Nq�àŕ'��5��5TxЗ��O��~�Fb�,�$~jRι@��5�##���"���li/�gz�3�MĠ���9ʓ@a�V���F�OG� о���3C������y����-�
B��}j_Yק�Q�*u�{�-����[-̯1��m=��Q��ߡ��@��Uv�R��۔�Os2�P�G/
��\�y\�����]#,�Q���gY�+^��Q���,�l��њ�OTok������d�D�t�!�괾�2�XlL9���M�X12���r��<�^�%-��]Q��}K��������
�B5���}|T� Yv��jǒ¼�:>"q��z�U�j�G�ی��L�⫹( �c�R�hyU_��J������1Qѻ`@kM��b}�4?�aY����sr�Ɔ��?-��s�I�	V"�"��$��=�5#�4�]�q.��1i7�Y��M�hى��ބm���_z�A=��4��H���OH�zl!hB�(�;A(+�����Z�{�C nMS�_��#��ᡸ�3�x)���G(�s1dBօu�O����T��:��ds���M/ŵ����5ᵪ����|B8r�}>Q�ew�/���'@�]O�y��Q�B/����Q���6�o����Qv��
%�RN�b�sVݾ����� �y��M\
2p�}�He����__H����f�f��;E��Ͽ{Z��v�͉qs��8�V����D/Ovx�a7wV���.��Ԧ��a��-�}yg���
�ݵ�-��2����D��i%-���v���g*>�F���_�����s���3���ʢ�ɷ�`�pv4O�cx�$�6Fl������>1{,��{6�$	�u��=Ͱ+S~Y	Oڻu�qp�ߜ%n�9���![η�]:�b렗�5��������Xhf%�{����c���
Rxj�n�̓��v,D��;/���Џ����t+�e��{�y�byt� �z/�A�ty� �䡑Ur}��U
�|��c%�P/$��%�Q�j���̑B	�%T�ۄ��Z�
�b֘K��.�����5�#�g���7��1�w
�^�KU��6&�x����_ĄXĆH�# n�GE��@/l���S)�v��ᘌ\�F:�N�׃��i'9�����~P1�0NF�`�~:ࡼ���EN��iW2�]���BG�_8D'sAG�¾\ykt���8\u�0*^N	�����NMr=E�£�*�Т�G�^s�_ªz4�ԓO<U���b`F��D9Z<*"f���H��&�!p�-��WT��ʠ���w���vV�l��|HF#���h�3�9��?���ߥt��R�u��߃ѷLUtz�Ch1�g�6\L	����p>tE��^�6 �Z��v;�Ԩ�(�y���@�%B�������E>$��6��q'п~�����9�a<�B����)ܜ��e�p<�`��I0�ru��}-���C�}#�-#�N-���%{�(6W�ތ<��Fb
x�Μ�ܸ�/�]�>v�7�L�f��+����YK����p�@e���IhT'v�k-7|���FUOن��F��tPBM{�}��(ﴟ7e��I��LM��@	2��2�i'S��Q�=��e`����fb<KʉUsu!��:K����	`V�FJչADVd�l ��s*�H��*����-��q�G��%�O��e"l=�����U4V�p��� ��Υ����Q��Z�˳.#����q�)�h�Nx��6��@T��00N��?o7G��oh�<w�9��j��є�/z- �����Ӯ^gt�P3�🆏Ȃ��]��dhܘ'k ����1��p����#R�� �ۊ��n\!���M���y��w&�]���`��Z�.U��x�)����]m�{��=<�I��j�B��o�I�L�O�߉��j0�Q鷨��q�/_q��Dg�8��V8�vV3�Ҿ ��y[�^����(��
.xy�x�炼��h5������,�|�oee�p�ԫ�Ħ��c�d
�nd��΁�be���$��J͜�+�%�_��w�"卬Q�%X�`�MnJs&�z�qmr���Lp�$!)d=�h�B�p^ֱ�������n�)����м��:����r���ފH���Y���<.�C��4�>�&̆��D�"��ńś� ����S�U�x.�@r�诪n�^J,�i���9�a�#��Z�Z�$����-TՈk�c
��j^|�#]e!%�Q!���b�ٮ����L�Gp�G-�)<���)��J����;�֘�j�Rg�^ݫ��������g9���=V�S�C����YhJ��O��\)M�о����*�Fb���]��wo]�9 �Q�=(�F[9͎��Nn�kyhT�WDN9��~?h�iI�'�MzшV�<��MA ђ�����/ɞ��EN���ַ��;r�4�z9O6��:��
@p_���4��� `罃`�3a!4|��A�-`m�BG��E�]z&ؖ���
!���m>S�Or^U�h�h����R�~&�/ "����>�{��y͞��S80q"z_o�.鏷��_(��sѱ?,J�B9��'��݄x8��i����[��/u!�.x�/T ͆�IFMr8������s7A�8<U�