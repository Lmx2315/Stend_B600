XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����R1B �x�MƘ�
m�!繒�v�ހ�E��;�hU���M�F,(��hI\��ة�6%�E'!�נEG�Te۾�*�%^mĺ2����d��Y7�� g�$>�����t�<Z�&�� �b�\�R�H��Z:�4îZ�2��j�&��6S��؅,s���a��Z?79�ۍ�0��T<M$,�I����)����vF?�j]�צ������b�+��A���^��:�H�S�Td�RH�]^z*<�c�����cH"O�����9�#��t�*T��Y]~����3�p$i��8sk��N~�Yw��v0�n�{�S��)���Ճ�wBܢc�Р��W_g��*ږ�Iys��ֻo{[������p�rV3�HD�[�O������f����RA�Kiy�T�u�k�V���r ��WZ�?�Y�hf�{[�'��Dt	�M!{�$�I%],u}ɾG�7��0TG ��N+]�J���,��y��[��>����
��y��J9�5qH��"�Y:q�5�8�l��رQ$u�������,f��J��E>a���?�ck4��S��t
C
������Bn��:$��f�$j&a0�KE@ϓ�*�V�@ݜV�ȋc��SSn��u�Bq�q�»!��c��!�Y;�3�]�H8�7`��{{q�][G��A
ք�hxV�[�� 'C�?��7�������,+��k��V�O���P� BZV%����K��y>%�+և?��+܄oy��*���cf�ߞ2XlxVHYEB    500d     be0���n��|:��0�����v �)��D���{T<"^�7֐�U/�\{�8z�G��N���p�4��M���qF��" S�ߺ�*"��/p/X�c0~��'-�OX̉�2�NxQBf�i�5~۴3���⫁����fr2��,�fL��K�Y�['4s������dA��z��7�<�	�`�.�ߢ��eO=R1�U�+	C�<��~�$R&����=7T�����v�fw*��7E�BƷ�&��*�HBi�\tl�v2>��emdD���iO�o-Վ?�)ɬ�6K�O05�u��,g��`��.��[���?�y�|���y��*Uq�[g�/�?��gL�P͞���{�YՔ ��} ������f鿟�%����v�7�r�\f�7�s�n����]�����Y�[���@�A$	��rm�8�HD4�%���r�dy�O�D�ber7�=��fBOk�?��w�k}w��h���*{?���aD����|mr�B: �TQ@�i}�C1�*l���BO���
�e�t����.:mb�]=���''�:�H=�A�������uⒼ]�����M�_�ʨ�����bds�'>�^��3�H|L�Rh�r@�`Ǵ2
���	�D�rUq�e���+`;���x�����7��������'f����ҁ����LOӻa�����	�w��(]�Pۻt�E��I���ɒ������OTX�[i[zQ*8F�`�:��I�u+:�u�bb�dR�'�i�,b2x�0�djNǵysY�46R�nCY��Q������-!f~;[&�_��c�fgm��)y��`p�Q�S���,[R�=Z�*�`��ۙ5C�/qj�Ma��:�𢽹�j��ꩮ�kؕ���E)��8%���AD�8Y?�L�#��j�vl1vO�TB"���
u��R_���*Y Yh��˶\��I\����\��A*��H�)c�^$,�'�dn�E΍ρz�E1�D����h�?9_h�25����>������0Q|(o`DF{7kqk�_�����O�GU�_�A�Z���$���8�E���kN���z��[�k������
m�]���:k���&�����-Y�n���5)����_�(����9=-O�9�����b����Y΢bp��Ta�3Ց��X�)sG 4�rl��w����4�;���4��va�k��H�2��_Pܕ@�el0 a�Α3�<��U#�A��"�do�*��_3Όok��"�Gb�$�)k�C�Q��R٩jKM�p���6ޕ��L���#�m�^~Rr�ÿ:�
�X�g�Q�?K��-�^�H��h�9*��\��/�"K����B9=u�p��8Y���[3ٍ�^��;��짒�X����2^�.�	�O��/�
9��̕��)}G �W�D%k7.��L��|X���e�V՞������%Oh�q&p�E]&|	am�� ����a:�
�hx��W�R2�,�tF�Ͻ�^�%����t���hk�PoH�{�_���E?#���t,A�C�EOc�>Q?�#��Oiw��-��Ųa��GT�ƣ�-�;f�T(�2�ˏI(2���5��� /�=m_��y)	�b�#��g0_"��jMk.�Y�g��E�������
ʳ\�0=��N�
l�9�eE��θtK;�<t�B�)ø� o=o�5����9�p�#Kl�#6���wA�g��H�<��0�]�(z3�?�-��R��,��B51�I�c����6�a6q5w���Ev	n��41b����%[�RO������KdKC���;��%
|m�,]���#�!oYSA>�ԧ�!ɐ�h�jMPU�_��9UxQL��,��x����b'/?�п�Љi�5qU�����k �x~���������$2o�j������zD{����)��5^�L�Sf�N{s4P��+m䇙��6g����D|ǵ(S�d����Z�i��db	�`鼘26i]�t�:��=B�6���w<��D3F���n��7GJ�AZA$ݣg�B<�d#��V&Z��z2&Qs�� �A���
15�������(�:;��e���#N>>wK��WoOŠs�J�����?��[��ΊY�)�Q�̂��A�q���cBu�I5`C?n�*o�_�;iǚ�㩬F4���*R�>:���~���`��DF�V���NV֓��\��i�[-��R_�o�0P��bF������ˉws%�i:��)#�ぬ�u��n<8VBߑ�ӌ�hP@MlMD��Y,*$��E��MX4����~6yP���-����Z�푮�֖l�oz��Gh����-��]OF��l�́�kD�5|��j�+�����kt��J����Y�����{��񘱪F��K����xcW�!��ԛ��O������ �����r�)9�!���8h[�v1���Db�v�-;T��h1�2c�Ld��(�i?ʞ?)�6�b:�rȘs��R5�tu���<�AO��b���o�8{�H/��TJ
벯< G��j���e�Za�ΨS���kXQ�ס�!�1;H���E?N8��5S�Q�Z���G�Ϣc�j�, N�l�`,��S��k�.�š��udש2)���~i6Ih��p�xя�IIv_��01��5��)ؔ{���WjR��/�/ވ�ZKJ��� �[0���ѯ�F�� ��Y!r��X<[�A�97�h�#Unh��hh, ��L�:��̔�0������Y�����q��q#��<��A�
�t�8��E��>R�l�,��!p�I<B��D�Gt�Rb#%r+�y���-���c�+���s�>ӏFUaAO���;X'�G�sZZ���߿w[ ��#�A\��6 ��ſ���[*���߱���j����;VX�`z��-�E�B�țQ�1L�H٢�$W�b�ga����B���)�����nI\��ӯ�X��8�ٞ�]�7����rⴀ[�0�Y��6�