XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��n�I=�=����K�S�|�p�>0�����yU�RT-6��Y�� L-�V�4*�v�*p�G^~�us�<v����%��e�t8�Y�E;Ʀ{����� �e�iw{.��4d
[�G��n�.I�+��hY��>وȕ����C.ǜ	F ���f��?��X"y��Ŧ�v6=�-���eW}󒄩N�߉�l��W�sc��b GثY�0q/.u���:sF�ղ��^�d8��C�z��P�B�B���R1�^�S��ʖn,'�$y~x���/B\c$��DK�7�].�`������+�j����m"��س�щf�`��?E�ghUO���]x����������� �[�E���a�n84h�-��>�z��R'N��'��@�<�8��Y����:_�(��5.�l�u�t�Z74�Y1���y�K[� ��Rv�M��d6��E}�|�!L�i䯷��cx�ר�މ�O�z�j���;Y�ZWB5������k���n�JI9��Y�5���,y���d]�P�j���C-�����d��D��e���6T0�$�W�2�����wO�JG��N����*zo!x�W(�.j1X�:w?� �N��o�=�<)�B���mmtsڊM�EmY��n��?���������E��X�N�e��Ԛ�P ���kd��l�����U'�?¥3��|�;��\��p�V�P-�To����}G���rT8�%cHy+L�&�o E��� �C>�y�%���[B�@�^�u6;��XlxVHYEB    1d51     7b0���t"� %����D�����|��	q,龎�5b��(x���%��E��(C���z���X���F����*�Cc,"����5eE�,���K=���ӽ����˰bg���C̥�54���Nߨ���L�N�&��V}�Qψ��v7z��ֶ�5�$��##�8� �]��
R#M�����I�GWr�{.�`���<:��'X	lLQcd�tUB�1[�J)�r,�	p؍�[��Am��Y�hJk"�ۼ/A��둻p���bmUpԑ��B0|��}�5T6K��>S���p��*쯓���E2Z8�^�Gt�1��"?Ǭ�7��<�:b�_&����_.�[ ��7�rYź�C`G��� ��چ�)�^�D����O�Q�=�~mm �N�vi���m����K�WA~����G�`H�{�AAf>L=��V�p1fRj�e~�.����>�J��5�9%��&�3���O6�����	��(U�TN)%Sֿ�+��,j�����_��,������y� '���q�kpU)I�u�XM�E?5��3��F\P��Y�pQ�Hǉ�7@�Ȱ+�e�ĺ��@HL_]Q��� ��βa�'�M��� �-�����p}�qJT�6׊�x���`5�$T?С�"���c�C�Y\IuW�M�����<hW�Ǔaՙ��ҩ�R��t��/l^"G�؀'2ے74٫s���4L�GfAڶ0���]g�Ŋ�����SGP���C0�g�Vz%&��C�Y�%h�V�Ҍgd+3nXcy����3)�Q�ͮ�lW}9C2�@~i믡?�,@�vޤ}iEn0TPZ'..W];M�S�C{I���d�v��YŜ+��ȓNόe^vo�aWJ�17S+~}XnH�4z���/�o�'º܎m��?��U�����IM8e"�����ZZp8ش.��p��e{0*�֥��/o�?�h>��0���w�<O�0!�{��kd]�:;:݃�/��j"�$Q�q]�}�!*i&4��=k��ņ�C��^@.MP;���KW:#��/��bg0�����hi7�P�].&���)o*��8�5<S�W]f4�52�o1L��#�ÛCWI�>�g�� ���E��$y.Ů��ud~�exQ5D��M(m9�s��b�O�/�>�"W1?�Ay8���[_���� ���+z��	uږ7�=�4�E8{��,۠�o:�0Y��SM�ⴰ�j#�ŉ"�B��bs�x����q峗���l�W��� [�2�Ӓ�p#&�ہ;���Szp^��=-�����7�u���K�����ýwŎ�rt�I�h>!�F����� ����+��OT�T�d�zk�L��$8�n�z-��}v����>�NpGw�}W���P�9n2!���P��%�frW�OP�N�}g�����������D�>�m%����`��87�:RU��oX=}�i��3�^f������d�X��"�dK�0{�<fd�)4{~Q��i!���0����[jd�i�H�*?1���I\�a��]���#�Tms$�y�y���G`v��D�,���F �|%"G��P�g, ��kY�<����M-i/��w����M��J��x�`.b�����W
Ԁ?��Xz�)֪���dSyx��@c.�b�N8��V|�Ѯ�qc����c���|��-�vC=��vp�lk�Г��s�=���W�ǔ�U���g�Y�K,�VmS��{X{Xȩ7�N΍�@>�(8�y(>Z/�Ԭ�kɶ��,h�I����J�K�[ȡS�Hx��ҋ~�C|�U��h́���>O�x0h|Α(4F������F����aڊ��K�.3��D�k��]��۩d����wݜ�|���8�K�ݺ!��&�i��Yr��|�|��3�G�]�z�m�� �X�#��f��C��C�Ě�[����u���|:�b� =Ovf����� ��