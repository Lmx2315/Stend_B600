XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��]i+!��Cge���J���:v��+���fR�(��߃���mHr���da_�ۢ��R��xG+ѽ�@Vk�sA����#!&��`�/��-�	����P;���/{~��I��c��8�$af�Lϱ��V�<�`����+@��o��S�ïu�Y��{���_T۟h`ˬ"�G���T�:�Q-ٯ�����Q6�ӝ�̓'u^�y~��;+�?��nWދ��4c�l/���h�]�S)#θF�Q�[A���i �r���xL��.��p���G_��-*�@Lez�=|��lS���.����`�RIiz���u�ҽ�(�v�w��[�]��g�Ϯ3�z#?�� �;�]A����!�m�AQ 7���0�=��a���t�(]�-\�	��+50�;���7�1wGS��2��v�@x�V�	Z���VG�?3G�kw�����W��偲���k>�T˅���2D��>�N�-q�<1�<�%'��gFm��8��~tU�{j�*8����>�&Z�Z_��F��ƺ��&��ґ=\��#C<,���c �uD���1�i��w����X8��ӭ�k�a�T�z�H�Ҽ8rJ�hjc8�h��pO���}�݋'���n`Կ�_[��#�Ӻ�������d�~�/�r�ɢ��+%6���b���M.%��7w_��WO1��Q6��	jO�x�beE�rpuٯ��K�̂+	����4О)c�B���=Lb��gox��XlxVHYEB    fa00    19d0�B�(&ÛU�/�*�e W� ��J�������!�uh���y�F��"�p�.��� ϴ�8��[ʵ����*( R��^+cm��WR���Z1�{#�F�@3,��p,�l�� Mҗɏsn]�1gشśM=��/ў�m�ST�#3_{�K�0 �$[���|[�=��Q7Ɯ>F��i?�k�:�8a,M��eg�JW9��������,
!�{I'}1�cr��O��B�U��/�qi?�h����]r�7��J�p����ێ
minmUY�*�������iX4}%�����_c�)���&'����Ĩ�l��Ǹ�b�h��ʚ��ͱ���=��G�����O��`첱#^���8)5���=بj�W��`�Bs�T����j�jw�\�=H2��V�W>�:���z]���L&�%h�j�a�#�s
�u2��6��M�+��c'Z�I
�o0G`��q��Sd�����r�lB�pxCAT`�w���7Q��h
���h*3�o<��>��./JQ"a�g
ļ�]�˚eNTQ3>��K�U��+�O�_}G�arB��Z�a��g���L���:��|a��3Ҋ'(�c���)�
cy5q����,;Ʃ�� U�~�=��y�ag���w	HUV;�g�H8{��St�pc��
Fk"��-�D+�8�'z�E�W_�Z *]��t��w�	M��wӞ}WL��<�cz潮�r9W$�Ԧ��h^��3Lt-�:��;��Õ5m�`�*��L�PTPs��a{5y��i#�ɧ�"zx��2��t�#�s�w7�Mk��)���޶����O�Uv��Bnr�`�1���V�N�M,�����/u-�.m�ɥ�����lNiD��Z<?�}Zw
�/_�@rZ^Żz��<��wy�B�����!�,��1#�Z1���z~�b��
/�b��q�m������$L��)��{�	��b�{p���U��$���-L)�?Z���|C�%<�xZ|~�R�P��Ǉ�4GtW�t��Dsn�Ǌ_��M-�_��Y�� �1+�W׍C�"r~��z ��&����%~��$-�-��A���2����皤�3iؐ��׍�v�\�er�3q�^r�H"�f�I'�x�u�D��@��F�Y��	G\�݊9�\�Ȳ ��&�*k:�ph�^ҁ_��<6mg�sq�v��s0c�[���R��Gw�&��!��r��E&3�4 ��#���Y^;3�?���J���k�<j7��@2%D�BЕiD�.� �\�1E��Y�,q6X�j"��$��_æ�(��MT�g@b~Ч��ȇ�F��Ef56�,���7MLp��#PJ�է!�5�
{g=�Zԑ�l�1� f
�#�Y)sf�m���"Pl�����������XU9�m���9�]1s"M)�K�5�!���75d�P���(��$$]�x@�Z �i蹸5Wb� ���}Bˌ��`�xʔ��Mdݛ�7�XM3i}�R��]�B�ԍ^���&l�9$s���ךP���"��@���s���ݲ�~�� �ں]��쁚���V/w�S��hS�"�V�N
�)��(e���!ƞ����1��2��ޙ�O8%u�V�zVD��e%e9Tщ�����_.��y�p�x]�� ��a���꿎��Ss�mː���_�X<��4���{1�=��2b�!41�[���=eʰ(�PO�����4C�ɻ�����mQ�]#�ȡ�*
�O��!��9|��S��'P_�aJ��8��������s��η�Q8���dyX�U�J4�
��A��EY��3���h3��3�����'��$v����k����o5DU&��
�E���}�N��u}]�?�d�\DlWg�:�)IP{iBs[%E	��f@֨���zWt�2���
?�]r�y��ex�h��դ��D��X���o3l�-l*�S�p�)�N����T�*CZۜc}V�!���Xw�V���x�a�REO]":��
��s��:L��	^�E�;�=�D�3Nl��A�	�")�ŷ�T�<�Ȣ��'��`��L����̤��}cuz<���� ����3�R/;�����Leev	�+D��_��x�����ڭ 3����	}V�d��ˈ!H������2� m��4�mz����Ϛ�B�
�9��kRF,�q�4������ZX�c�=7��=���(�W�vx������e�\|ѝ_�d �/3�<Y���I�1����&�?K�'�%�L0���/��dL<$;3�cb;�]���Ú/�����ۣK<Pcs@nk�^TL:Y~�����
���r�]ЉLǳ`�(Τc���j �"�!�#�\k���>	�Yc}��5 ��0S��X��vR �@�#�T�"'EC�N{�U2
XIwN׿�դ*Uz�ٟ�uz�Sq���92k��/F4�9��o��6u@�m�;��3gy7�h�3�F���#5K������0^�B��i:�P�9�Y�
���)�����:s�ޔs52�1�d:rQC���������5k����k� ��u+Bj��v]�?l�a	H�p���^k����*���L�fୀIŋ��Iik5��q�i ���g�h��˛)	��T3��!8%Jm�?�0�B(�h��+t'Z��g�)�"��^��
�������p�mVt�$�8iL��\@���T�2��/�Ͽ�,�\޺ү�]Vn�&�����FJN965<���&��K�|��݋���(ͩ� T����u�{�J�\![�	���Yd�G2���N��o���,N�a���٨3�k�n�M��*LГ�ԫ�@ø�(3ǭ*ةO��e�9���D.bH���&컰①U�2K�Je$@sK^����Zq��L�t !*�nMUw?:g��Nw�7W�2L���RLhf�L"c�����
��A��m�_��(2Ƌ��綥��W��%��oO��BOr�1i.V�z1���"�o�F����]�2�!����k��Ι'hqWVs頚�^����քVe{��BZmӇ_'W�2&�⩊7��(κhwb��=p�$&��	؍7?��]�-����)?^Tb$�N������_e~���������NI�6L�j>[OZg�y�h����톷�Lg�c�t)oF����)�6�lFk�|B3�3l�hA�$dUN<�TP;�@y)��v����zq�����N��,�|�k�=N�P\�M�ڄҒwU����n��sEL���x�}�����׍�53�sV�H�,��p�9`��/b)^R޴����1��,C����b��*-gB�b��Ga^�� p�s=˴�YIg'�)=L�q�/VʱnvHV���,�;}|��iU�II�6�|Ǆ�e�eE��]��6rit���Ӗ�&��o|[u���_��j�;��F�i'��ʬ'_u�{�f�\�����m�j����G�C7��V���)��ӗL�m�;x��T��k�K�K�
����f��%{RT�;�a���wQIo"U�����s5s���Z���p��B`qTH��?���@dW�J��"	��P[�e��~��x�,&�˕/NAz���>�Z#(l`h����w�a�ԪB�)D�m��h厳��$	ckq��4
����a%P/K���������=��P��X
4cuX5A`��^���c%���u����\��_p�����(݊�2i5"^��JJk��ܞ[TBQ��(05ʆ��n<�����	�J�l���Ҵ5���ֺ�M2��Aũs���J���c���׹�#8)QS(Xm��	i�G��oR�Etü]�6	E�E)�~E\�[����Y]�=�4yL��~îy�bP�8֓�x��вJ�T�A�6�K�i��w;uq蹾]�ëKk=Ŵ��Z��8�pF����5�&Ǐ�ޯ� �9&\"�~����K6=,R��9	Ȼ��~3�����N*���|��x(ëm�;ڲKqt�{��O^g���}l���jz�ß;�%��	��}�BEy�L��w�^�"/�.4J{iz�,�+���KԹ��(�Rw�b�Ĝ^j ΐ	��y�?XpY���U�}J���lH�~�����2�@��Y���݃"��ꌒ�?H2G�leX!���䤶�B�EV��8�����B��%��I�[����ed�����-횹J{��⁉X�	���c
]�'��*yҞ���Y4ھ�m��Օ�빉k3�Ֆ��|/��U*�!�rAW���T����q�!�"# 5�����b�ϱT�A�;� ��R��"V���Y��>ᚎ�F����Z�9�S��`|����-P�:e�έۦW�l'Mw<x� �/���s.�t��FA���	:��s��X[��Y�8d	,�E�F�'p���.�R謇BA<b����"v)�9+
��#�7���g:��"���D��;��i��w��!�*��J�O����L���f�o�=� S��ѓ�|ƽ]���@�T�wE����s&�TDoپA⥱�umg~1����c/�)@{fӘ��-��j�>��(��~�-㭱���`��5�2�n`�3���Y���q�>��T����G��A,J�_H�S���b%浨Hɳ�M�D�px!�����ץ�t1��\X�/uc�Edw�J�' �G	�,?�K��i��V[Iծ�br%��eE�n��j
������������2��(E�_�#�Y���,w��q�]%n���A���S-�0%�MۚV4mRj����B��˄c?���ȹ@n���;�g�
c�x~�Wk��z��A;��ﱮ��O:7���-�L�e7��V�Pe�!o/����{]�C�!�B�����h�EI/d9����Df�F���Y��E�o��;��+�?MƩ"qP0r
g��F�����8ض��E�y�hǬ�\���8ZKX�V�Э�J�,}2>�Ìe�Ҫ9L�`��u�����j �\��L���D��xR�$�eM��x	��$���&겺.���]�߈�Zw�4���/k6���fݮtN��1�/a.�2yIۏ������Vf����iq��k�z�ۓ�3����Є�.�_����b�!b���-�y��$U�L3����r�����*w�����'ۃ7+��2�g!no�|�Si����>
�c2�cR�9FЍ����0���q�'sn ?�̀�����{Ʀ�u������O=S�3~�>/�m~���)W��(��O1�����etv�̣�4�&���Ğ��0�Qr&�ڣE1�;A��,���p%R�5�WK�y��� T�X�8��2tCp#��%�@����;�U����ZI��*�qj���8bI#&�2Z �z{�=>�
��|�z[�'��AX�#d�x��: ����A���71��6!����kO�'�ᯐ�M�L{ܯڳ��_~�
����sJg�o6��1�[���2+8?FN�;��T�G�7�K�L���&0&��q��FsNw��n�.0��eA�-7��L�Vd�"j��?�$p��	�ޫK���Q5��U�'��g�r�*��O&�E�i�����bl}��mx����z�9Y�U| ��Y;����H��k�b���J��1oJ�|�riy��]ms�e���Ǣ��ed����aFWf�}eEbH-��p،��M +p��lHo��pXe���&�V\�� �a��<���Ch#��6XW(l� o��)sK_�.�C��9��Q�W�Au���Z��A�.��!�gS;h<��)s�x}�/�O2����>!F�ggn��7x�pQ8&���J0���R�rƽf�����V�#HD�z͹bl\�,]�eIޢ�n�W��B�p���1c3dJ�G��SD���d+�Z�rO�1Qv�ؑ�����Su�����]m«Rn?��z ��TZ?M�N^��n���V.�!{_ K:Fm�Dy��ƶ�fGQ��E�'�c�ʃ��$���5Ȯ�95�$M�6c┅.��";Y�����\$�Ӿb><�~q(�3���Gq/r�8HOu�JB��a^�ȍ����R�#�����9�2�|:�/���)[g�ex�l���Wl.�B,���%r�U��'N�Lo��>/9뿟������{9?!.���ex�C��K&/B�ھ�բ�-`�tė�,��ʥU���&B@�%|�2��ꠂ�po9���Գ.��SyCB�/f	��E��dF!�ʋ�˧D��x��EHkj��s���6��y���h6�"5��I��nF�>�_��U��(�#�ŧ�/>b$�j�W�ZaN���18x�f��ĩ��5����ޯ׼��a�Q0�7�$ع�	M��TF��i<��E���
C���<j:O���JM�����4��¸�@� �?�����c?i~QSFRȚ���$*���}t�����FE�=��B����yF߇��=�֊�6?XlxVHYEB    fa00    1630��p\�>���w&�� ����C���۸��5��x����ߣbs\���H�+8�U�a�&юWd���tM���o^G�z�,�����JA�z�?ҏ�wn�$7��`�=čp��_k�6�zgCfx�M�k�4��	G�%bS�z�;�4q���dnַU�>>Ar�ùE��V�cٹ�e{���t��b�"�r+!I���z�S��=wt��~v�ʋ�W<됬��䟣1����9���n@~�fwH"}�bu�c4D���f���N��X�Igb�zf���A.]��$R�W�DAq��1�6�x��=|:1����-��W#�i�q�g�Y	�_U��pTϹ������󄾳C�&R�ئ1ޛ�"6�[RB`#��s�)8)�e�Nmsl`Vo�s����%J]Ïo�;u���T"�a?���;=)Bw��	�(�5T� U3��^ ����w�v0�kǸ�hÏ9��j���M��EY����/�ƞз�VQjF��q1�4��-�
�A%�Rq��p55�bX�� ��ȴO�mr"����e�*��[��B���ʄe��.�s��9{�3i�cu�v��&o{��{�~����6N�0e~O������D��9o[�N��9#���O�][~B=s�̡G���W�Qϻ�ҲN.�����S �w����vC�����8j4�tC����Y�n����.u�ص_8�:y�Bֶ����r]�d�J�TN���@���mN0�U�1�]�Y+��P31�UL`^�X���p���C�M�ߺxS�C���>J=����o&+�h���C�"y�'1̪�f�cN�uZ\�O;�O:�AP^솼�k��e�Q���"iڙ\�:�W�pI��gP����=��(�<ox���dحN�vLN�	�Z�����4�]�1Wz��(Ÿ�I���f�/��F�n�o(���9jƀO�Y:^
�����,l�]��:8�O��{�sK�W���r�K�Ah�(?�?�$�Iȟ,�1�����_hp�F��eDRMM��3h��'�� �R�.b���ӟ�X�X���E
�>ȏvPup�� j��F[�ĽY����BaȄ^�W}���I눕 �̎�0M�:՗8L*zvaTΰ���Z�Km�|�^�#lLؓIf��@�����uU��ѺC��$�S�ƕ]�!ݕ�bB!k���m��7be������.�T�|�T���N����1Y:�p�+7��<��J3+����U3!xF��!K��������w�c�X�
�Z-�/N'���v;�%���xu*��`;�������ZK#-N�O���K����oc�ʰ������pi��W�ݚ]�a��*z]�����'<۵(��/���k������c���i���%��#�z��k�YYĵ8P	�����4b��	�&��7�w��ܦ+�G�M�R�[QK���[ID�W�2+�[x�i�6��A�c�3�V$rm��vU�st�x�^P�u��!����ϖ-^��TB}08�����P
��b�X�ͅ�z��W@��ł�8.w�g��vI����+���eVPe<d�v��ٓ�
�!k�f��M�b�j��C����x5�������~AL
QR���|}���B>���PɊ��<�K����b�J����t_㓑��Q�	�:��\�\|��Q~Ye�v����K��^~"9Ĳf9�=j"8e�e�+���KI���H�v�BT��
MLַ�4?��>>˱��(v��G!�ks���
���"*�T	�Pc��k�(m�8�b5��D����P�-|ԡr�ً��R4���8����e�2�ie�?5���dp�C�C*o-�W,.���~�X��!Єw\$*�-�s��Z�n�i�+��B2�+�-=���@p�d�#_H�<�Sjx�&�>�p��lx3PY����~VwГ;	ڌ4f�E�(�fYU-���h(Mc�B��P��L��t�^ѫ��oA����yG��=E���魩v�������Qk��t�v�m�3�ڱ���D���Ri��r��-�'X�o�#�C`�E9�H�s�mc�z�ꎨ�)$B�Ra�t��=���T�=\�Ъ8�����C2 �2����b�4��e&��	�����=S�_�z��T#VU6��ć��P.Y![x
.��d֏���j^�s��	7�ݰ�^`��"��^�������;4��� cQ�Xef���_f2�6D=�EE�>�b���rP�)�Wϸ7�KA�e ���u�S�%� �̄p���l`��u�_�,�� Qh�>��f7�M���W��ԡ�^)|4���R<!�Ć0�*y k�^�2�|O���~W��`���^��5���ܬY� �ώ/���NH��w���d�ǩC4Nn=�~n�I/��%��e�f��Rx�K�A��L�NW#�lXkb��԰^�Xc:3
�o4\)!���c��&z(�+N��|���H��,�WB����߮N5�]ӿ-���=^)U����������kt��\0\1]�Gd¤g���+$>W;f�g�&��oz�g�1�F����d)/�	��%�5�&\f��$oN�7�HD���n�N��A�������)a�|��ױ+�|Y���*�e͛��M�X���G+Z^?B�u�$)�!%�x#��K|�ؑ�(�u�3 �Nɳ'u0�MHU�܏��]���{^s�"��5�����d
���đ�['R��q�8F��M0N��5����9�����-��Y�-�b
�lԘ��/����ܴ�{������I�.xK��������f�����s�4c��Z���`�Mޮ�Ĕ�G������`�� ��k���EU��P���z~��.+�[?� ���gZ{��z�/��I!�*�w�%�=9 w��Ƣ���۱��۔`Jp(�>�F0�1���g��ۚ
婫��9�����&]$ho�U�����l�ƒɰ,G'���M�!a�G��>��a\(�H�M�M8����r��,6`�~�N����8C�b�}��A;=��g�	�BY��<K��������'�Ҷ�����9Q'^��L�D�\�L9���e�����T`@��7���y�ɴ�D�3R�_�]�Q�"i�;���s�W���䣵zÜǗC��V��,�K�h���WS���^�%&#!݃і+�f�Nı}M���o6ݰE>�?	�vISu5�Oi��x!�P	B<��b��ٻ��5��1�h^�[[n�3e��ћ�M(����hn�����̶gߜ��`�m�x���ER��O���#D�A�[�^�W��枝���ɍv�쒠���ӏ����b������ϡ5r��N�ؘ�Z�QEƮ�ײ��F�^�{��k߸�h�Fxs[�3�Z���Wj/�YBgX��B
G�0q{���GQ����%�̸���@eqs��2�d�"�t��^~:	�4�?]�m��bЫ曇!
T�l��fl�RpS/~��s�aŇ6m�`��(�u�h�(!f	
qi���%���x]��T2�YF�ς����C�!ĹdU�2��3¿e�H��䫿X>�Bl��;Y�
����.t�WGGu7}��O��V/_��zC�:����`Sx"�G:]�m~�V���$�v��'���3`@/89:���Ǐg�L޺����E���^/���[�^c;CK�EIEd@�iu����z /�p�g�*%A���m�E�M�	O�-��WG�S��T�<O��������r�}kd��4�y���b���
2WR���}�'�C��7�b��1:��Q�#%�'��9���9'��^AC����=���'M��B�7�f�7F3mN_�}�/BT�����N�R���א����u���p�)�(z��G"\<���( pP�?~˒u�&�%;C����S��C)�w�U�>��0����7¼@������9�(�4*�_!$��a�zI� m�hݔ�ot=�(�1�:�uѮ3%|\Z\x���\(������i�W�_������*��c������@9�-5k�i�e��tq�*GT��`;5~�^[Ȯu��R.���߾�m�K4��ΰ��cMN�no4V]�Ӏp�V�VD�x���j��$\��#�u�u�;:7�C�eb�I$�Φ��hgǼ���zki�$r�8��԰R�Q�B��(����O(aD�Wi�ʅ����^)�cPO�/d#'���j����u'Brƞ�����jI(���[�X��������y׮vE����K�`4�V����&5�"��r�$�5�<.h&�+�
q�	��i!�#|v[=C��z6��i�hCtЇ��� 
��'H�( }�:=�~���U�e�й�����8���(W�w_�%�|t��í�֧j�Ђ[��#.���
5���>}���-�\���Y�+,]��:ƭ��\��/d���B�,�=�L�ad�ǒ��:�Z0̈́W�]��l�s��|	q���*x��a�Q�ٞf b	8���{�����l��y����yf3����_��7 �o��Vs���q�h��0��1��b�4��� �oi����s��3m��^sD<mNI�	0��;�YZ#���L��q��y� ���g��қ;�W+����3
�f;�Ib��@KV��ZP-��r8��>��{/L���o�qƹ���-f"�?۵�"��n�»|vr�=�v;�{ǸՈs�r���k��U�1�0N5�G�����-��N8E�t9�ē�"�����Q�fL*JQ�k���w�Of�ΐh��R�]7L�NʬT����'�I��Y��i�'dS��=�n5*�@	ږ؛��^�b�b�z�Ζ���\�zKb�em��z�'N�w�[�_���&��#yE&V��(Vޞȣ�|�x��;'��Dӭc`!��09��)ͻ�f�P�#�w��X�����z��t�*���,���KG�!ȭp�'Ϲ`y� 4�e�}!%�턐���=z�~�H��8�\*[T��J�x���;�7K�H4����z�5
�Zm��Y�jؔ��5������M�'|s;�)ֽ�|Q`�� ���ۧ�h+�������ʶ�^��� t���lm�0�~�O���T߰kV�
������`	/_p�y(3�����v�-��d����
��r�>k#��e�p�$PhFS��rr�ߵ��` 閌����?_J�D�T�5��ܪb[O#,��4vM��W�V�F����4�̙�g�q���+�W=NM�Jsl���;�ŀ�P�dZ�^Wp�"�q`��gY��f�����&�H�i��!��z�3��4���'��N
�|'D��{-��F�������׷[�]�do/��Uk8��HP�3���Ljva��Ψ��c�����׍`�ڄ��.V�y2��|m�X^��f�O�ϛBH!Bѡ���F�x��+%l���,�<M �N�_WW"�)��s�8���$�<_��[�B��2Z�5��*ٝ���̼�X���|��W а���F�sv�GW�ڸ��Zu1(�=(N	H-`�T��1)��4|�]:�n��9�U!#��]}�>//��;�˓�XlxVHYEB    fa00    16a0��>��VY�=����f<�t�*q�9�����/�+�q���%@>Ϯ�P��j*��V������\)iW��ZE�e:r	t���ɤ���̃,��������3�uE��5Ԃ�,�{e<�� �8Cl)21N�s=��GOI�(�ݘ��:�!J��zà����� �t$��2�����5]�J�"��7H�� wA�����5b��س���T���2��l����|�
����X� *���W��4�����ݦ��O4���"�P�2�N��?W��]�q��p��� �ҽ���׻�1�Ć"�mx�:���m���C4���@�2;Jl����O������5��
k�6J��d��(���8�:��4M��cx-^D��@�-��)`�-3vY��,���IɰN�ER�'N�ȩY��r`�XGLIsZ`}������m��ʛ��~�jUJ8�(N��>8�{� �F�Z"I�y�*m���_�Pc������=�A0���Y�J��j���n8c9?�q<o�0�衇3��*I�C��v���36�v��_~w�OR�6w�L��%���� Ǿ��^a�^���\Y�F#1yl_�<g��qV��O)��[��\���}���se���Hf8��qN/~	y�Kk\}�3��t��O����t�����n�>��*lLm�v?�H��`69u��hTd �8Gx�./ ��8���P�e�nf^���7��u�v`���D"��;�w�u��2��-,$�q��'�w���E��c����Wl�,�?P���]?�+*����n
��Wܕ�A�V)A��q���pj4}�ʓ6+H�8�u6���q��`%Ҏ��pf�c�O% �ޒ�_��
o1$6��]r���=�����C(Nұ	��c�������{C�CF;�ˈ;~�399�����?�k?�3�"���I�q�tSYfV����:%�[*ePa-oi
�u��,ŋ��5���V�녃���5��	�S����]"|�8�
-�w�h͠�:E��d˘/���@���,�:A�T�s)�����"oi�B�)��0��EoH�!���B�aP�*^QC\�	 _�X$ph�9�8��ϊ���Y����=��-�8��6]�8��.(9={���O���X}�N�D�d�Y���#-�mXz�P��m�R¦Q�><�B�C^���6��0���ؚE^�\��km����a��d�F��!LN�W�\�{�F(���������.ݍw�F-�inV��iu��~����>l΅����Ɠ��-���x�?zr=
�j���L�&���������Ļ������`�D�RP��$y�*^��J�I�\`@m��
�?c�dA�i"��<����%��"J0>N���q<[�f��Z�]o�q�ǁ���)H�7U^q%��ăd?��]�)[~�!F��{[�1��wÛ���]����Ɓ��(��_�X}Q��^8�[Du���!�����;�w*h��a4��3A6X?U�Я��.��J�l�vJ$����(BG)~�=���yg��y��'MH္2^�B���;q����(�@��%�U	�B�G���z��#�$tk�d�_Qo�p��$��N q���^[�V\ 9~N���B�3��n�n���A��"7`D�zP��AWy���k�0�%��k����m�$H�o����9)5|c�K�`�o-��"/Q�C/�z&�嫭�t�'E�Zm�h�afo�<�F��\4� �jz���&KJ�xM�W�kٰ��"&B�p��F(�1�Tٔ�~~%��C/ܔ%�����d-�#n��x���Rak��݈�����)]�:���x���*��D�^V�-�8R �ܤ�¨�1���}�T�g�n���Z@x���-�g֛j�n���+w��[���^5R��p�w�"%"�?,�e젖�`W�B��ЙvJZC��\���~/#���,���&xЙt����m�8[�34F)���r��d �(^�& ��25k�4T���{Ixu�����.�[% ]���s��*�����
7��h���b�t��UT%����٬m��| ����p��BW�W�L��C�p��0K�i�d�ˆ��[���S6��rإm��*�4 LAl��*�Md����ZT��ď��E��z-���Uȭ�������/����;�-şN�{�盟�m��Y#��Ke���WJ,�{ �!|���<�V�zє�q�!Cb1]��YRg�򣇷}�yf�(�� F@�-T��S�H��\�%�텀�P��"��|���U��t_\�LOf�
����5�.�W�U,�2�F'�bCl������h�!��2���y��[U�B�y���TGY��_��+���ĜF**�[��Z�x��x^�k��Yj<r��MK���ҟZvam�&q��w\��	�E��V��p��d�@���������2*��8�' 8��8�*DY��U�0�5w�!v�.v>�+����\������Q/ī#o�3�N!��R���)���D�:_�W�H6t-}E���r#���]�p����B~���c�S �f���yR45�쒊y/�ӟBӇ��%���0�����ߪ��^������Ӭ�_|�{� EJ���nsI#A�vQ�5y��W������b$]��G7k�)�,� �u
�T\�b��L�i��*ΆtWFe�{�N/֨� :�=O�$x}�zxHY�*ݡۚ����W��-��q&/D�s�˛h��j�ύ���oN����ܯ{a�>w���5���HcX5�r�����w`4�^� �S�@D3�M1s�x�"ω;$���gK(ʫn�.��Um�'6�ك.g���f�YԼy/P�>~k*��?� ����sb�տ��&��v�R�@��7_>D�KB����5l����Ov�D��_�*��m۱)�(y'���ߧA%�YD��`5 c��M:�9HJ����'�2�Onlhz)[���$�� '���yk#uEyYRv-v�@@��7		{4�F^�J�~n՟���Y�K��|xXŢr�g���;t`�����OV?���)��LB�z�fё�I&*�y�Y���ae��S�Ly�S���p�<�����w�R?�3�$ �mhJ>���52�1�sh(X����T)�E�0:F�A0�v�dY�������*�QD��@��w����&�y�R��6��D�]nɥ0��������#|�m=�eՑ��yY��x��7A^�aB�Dq��&Y��i���';�u��a���ڠ���xEJ��Й�̰�sw�U��K�-������eV�9.�C����YwhD��7M����syKR�=�5�/��9Y�d�2ܻar�y�.Q�\��K��3�u;�q��o, C����"[�=e�"'A~i�F��|��f�I�^�5X�믍��IģE���$ �s��4?z�+��#�� ����="�����Y��1}��OT͢����+��?`�Ѱ�$U�d�Ol��ݿAK�;G]uÔ��6ka�Ĕ��TG�!'���@��7��_�J*86�#�6�*�G�?�^���¹��FAg@��8@�E��V���r�&U��m<k� +8e��qGj����pڪ��D5��йM�w�'3?�r�	����f��̜����s��U�gc
}	G��}_��>>��ŧٺo��U�9��G~5fUL���������$z�u� !m�Dnݮ��X�I1�^�)Ra�.x<�J�P:��u׹�X�c6�k�=����`��Lt}|眂�_X��b�}�0�V>�~���Jny����ގ�F��L�T�VV��K���xiF��1<W�3XT��r=1-�f	�������.�$K®<����5�ڵDC����uI�����r(�g����R��bpC�`]�CF�T���j�d�&o�y]�H��Y.��WI�B
Xcm �!ݿ�eQ�=}?˺9�d��ss~���m�p�]H���-��R=t�5b�)�Qn����r�����@�tC���ސO�[���������3jD� ���AAg2�<� �b8%�B`O>� �a���bL��9w�YB^�E�̪�px7J��)D��V%�m���נ�6/�~�J���OF����
���R�h]}��,��S������1�&�j�)�g��rf/7��9����پ��`}'U�����m ��xz47)r˃f�%CA�����
�W���*&��F&}�@�s��C�*�p{�p|l��Q������U�3^���~J�����6�o�	^ʦ	�U4rw{�_xQ�p^� o��Jҥ&S��M���Q�Fg��TH�����s�I�k��u.f��0��{��%�~*��$o	1�r�E?�TI�j�,�aU�Xd(�7=M��5h���m ��y��eK[����:�!|*q[�#s�OTT�z����cU}�$�&��5�k:��ρK���|x�"Sb>�=�@�FT�b\���%����(��8��i��P�F �i��,��v�t�����	�)�>QΙ�w�8m*�	ij�[�0�w�T���K�-�Mꓡ�{�P��/�EĜ����:���V�I�T��sv;@qA4�����痨�C���]�Ѩ}+槦	�R[w���4vi��f�s�=rH�L��s��j�R'�_Ӊ9JŶ\���S�W��X�S��I�I3oK�ib-����nz=M�1�Jxߩ='�(=�?�|��,�P��_5e�f� "�����|��xϔ�߷{�Fӵ���C� 0Ğ����]���NH�m̒+�\A��k�ꜱu*���߂��'xС|��j����i}sI3,�!o0�"��8.?v ���u�Q�rW���̍��G9V��oq��"��j�P<���>����{�0TȂ���ɲ�M�c�ћ�Ocq꼒)�O���b��n����o�u�٦t?�����ƧyK����y̰T���@LeHs	��o>3����?�&9W�f��#�Dkk�;����m��Y+,�\����u�˫Rz�ܐtw�f���!y�D��;����,�siJ(��I�~l-4�<R���d�p�j$9�oқ63�������'�r� M1�-����}9��MBÓϴ��밝(��Y�o�ȫ飝��K��*�l�3)�r�K9Co�� XdG�{���B�
�%p�I�W�����*������}��ꐔUI��V�������A��_��ѓ?�'a�����!���exY��n�i�Sw[mq�S��Â����B<�����][9P|z�M%F�&,��n�� t���WH�X����hp�ˈ���D�#�	������c[ź��5Y�壁�g��L�d����Xs���U��^dnP����x�XcK~��B�X7�����`�ʨw�>��K�U=����+�An}n��a��v6�}�?La�$�F�����Ɠ�4��|�R�p*P�Ѫ�B�|
@�HO��l����_3�k��>G;ƽ��2O6+��L��<�hC���S�/T�M���U���p�R"1��Wӥ�2 K��<c���	�r��]���dz��*��,�r@f[|T��CXt��WuJ����Z&���"D�ԵI�݈��0F 8�j��H9��r�愱/|@�yl׬y	��]XlxVHYEB    2889     400z�+Jl|�P�V.w>�����\���n�x[fp���U|��r����8Ą
/�>ԃQ#l�::k/�&�g�'A���M-�ݔ���e���;��_u���qg���s����ԟ�FʠQ�u��L�RSIc�z�#�	�a��Ar�w��.%l����8[��0��	l�E�S�+�@��5z�i&�E�n:�#��A���ڟ���H��Q�GEeO��o�ʘ��3�ڲ@�^ÝyF�jf���Y���
{`B�_PU�K"D�^��D�]�5�!��Q�?I7{���j�a�o�&�B���[ (nFLi�=���6�T�FmD��9�����=��5jGװ���s��-�&)�Q!��l�Fk�U��������,�cw]_O�d!����+�EN���M^3˃�/�k�f(y�J��ᚱ�ڼ���~Y]�*�`��yԴ��\�H煸Zkud�L�Z>#1Q��[��kb/���(�7e��V]̥6ű�QY��z�2��Ż�']oV'��tP�k�a9	1�׷��(�vVu�¥(4,m͵��b1��v`��A4lf|��"w+�>a�(�B���^b�f��xZ̭��k���kˬY�H�_��h9��XXj���#T��t�����i䙐�ll�~����I��K
 c;Q��ڮ�g���h[��M[��rr̎��M"W���̦+�(@����*�GS�̝�5�}�cCT��YdA�!��ӣ<55r�;O�(�R�������A���X�E��M�X+��̫;����]����*v�i�@�0Ld�p+0#8}��Ұw)�`P_o����I<D5a�Y�6���+nX'�D�'�Orwպ7��U\E9� íD��~��:�^�7É�4�(�j�R ]|�����#x��9����v���
r'�V��������%�&���#�>�`t'���m2�IQJ�, �Xf�&O�f��
��Fa�`䒺~��ܢ�j[�csG�M�J���p�