XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��0�� sPQ�8�J�m�o��r�jWԋ�lM*Dt�C��Sکd��.z֤^���ɯ���~=��0� �v�v�����.����*�F�R��j�p�c1��al���t�P^#�r%��{7���,Ä?��l�$� �-��N4�^`$�Wᅳ8�Y{�p�o7�i������]~nJbLSc���'�j�c~�0�֎(�T8n�g�g����dWD��P,td�o��oI;4U�!��91V#�o ��2ݔ.߈�Ӊ��?���9%����]xh#h��H<~��Kn�,�l+L��[����R�z�4�?������r}��ڿ��	[vFbO[��q��-��:�/;�M�|\ёs�/'C�����fZ�;�	��.�dY�ޅJ6�`�m�=��hX�4��㎑�օ!��ᆾh�b�j�3~���'CV5�@��8���g�h�$%�,U*���Y� ��	-'g��"��/
+��?&I䈖�57�'��/��U='�)23�b�Q��R�d!>�&!5�!�Bp�i��x� ���@A;�GP��:�������:�3#�/�߄wv���8$��H#���_0�AS�������v����V~~;�𝫧�$�?z6�3�_qXۊz�U��Ա���x�9�8�+�S���������`�Y_\+J��=ynW���������2���r�f����Mw���(	����.%�B���'�ѭ��GՏ(u2�^��J��0XlxVHYEB    2b30     a30���i���"F�{�DtUT�:O[�Z�mr��U�0
�m��,\�� �d95Z�><8�t�G�X����Y��)0@�v��á��AAxEd���G��"���Te�t�n�J���L�a���X��6�����be7v�nhͬΖ��<(VdI)Sڲ=����y�)���ŋ�8-C�|�G9�M��p�➵jb��y�"^�4v:��yOM���H�@�<??mݑ��|b.1P�.�����E����"����:yX�N�'�U��@#3�TNB��mTU�g��RkL�d��2Uѱ��]}k���e���P�ǔ�(dE�7���;�	Q�y<F_��t鰪�k߄�`��H��̛l��,Hg����+Q0�ڀ�}�d�F��~�^cyT=���O��k�ɲ�v��഻�A�n�F�.s/��E��c�F.`V�D�!��ͧ���=��)�:2��5�V�XRL��A�ݣ�3��8��l9unb�Ԗ��g-�5��U҃ .�詒��פ�1�<�Bx�#*��B0�Rw��O�
$���U�����,��q�B�E���l��f���8|9 M'�'�Q>J
1�����_OPR�W��4g�ٲn�
��W�w4f�Ú�ˁ/��ӛ���]������!pR88j������%�����vs��^���U�K�s,m���l$��-]���mvk���FR�K���Y<��������N$,-�8�� -yv��@�����{����<@h����6�����.@�G�&����ѵ�Q��QjI�R��]7~��@����[o⮺�ې L��Z���gg���������z����arG&Ҽ$8����Y !�M:��f��e\Lm��~���������t�ǥ�����Y2Y{R�^��ݱ�j�Nْ�[
�S̩��v��1>(;0����`���5�:8���Mūtǂ.���'�	��B{iq;��UVu���M*/7�n���Z���v(��vl)�����H²�xp]�c�Q���e�tޖU50[!�+ʄ@)�H������{-S,_r��N�{�+������`NI_���wzH���9a�UPU]�x5����P��LùϘK�Ȼ���� �� >.�FY�Jk9��D��XP/�	j�^Ж�v>̜Kt��{/D}@T1������>=���Ə��ƃ��\�v��Ƅ�� n��BpO6�
~�}9DD����3g���D����^d�5��`��	EB8��t��D�J=%ҋ����$u%�>��n�Ӵ��x[|�d��2!��=�T�2Ϭ)��"��(�2\��H	��ۚD'ZMQ*�/�������v�_z������cL�d�V�y�ok+�!aM�?�Q��(k�cj^�D�n�L��r�@�c���1>�2�=R��qm���!'bu����;nL�f�^l�����z��]�q���R#Ƿ]�����(�3����#(|���c/M�(Ղ�{/�t
x@�>�[a�/v�e��2�sy�ٚx�\�5��g��2k���Βː�'+륇sp3�	/��y����P�9������p�����P�E�c���{�����@���T�6�emH�����ߔ�z���0mf��Á�Ľ�v~��N�+E@)������0�W�P�+7B��Dcp9I��L3�h�P�:ZW.8�ψ�t�u@EF�ۀN���Y�j�d�}}�8	�����I��ހc����L�1�����RZİ\Ȩ��v���A|M�h����� �F/ݽ|йT�t)��֠_��f����O��<���%-��X��t�ೂ
��=}�[̫)�j�ك�K!�l�}��t6td���C�1e�N�v�_69��X
���Q���A3�6�@U� ��%�r���D�(_����x�p���h��2m�ΏhڑJ��D",�2��|W�����qH�g)��A`�j�v��&��5(��/ &_�ײ�)[g�8���K|(�
�\2F7� ��B�࣎	1-�������gNse�d��&AF%���A��L�X�d�������	�,��<�C�o6_����>��#��swa�Y�
"�Ln�Vz������/Vd��<s�_t��JB�����9=�>�px>E����y��:�'���c����dM�Vy�{*}E��Z��	O��5E�~�k˩�� :��¶r���0!^���p�e�����LW�e����ү���Au�$t����@��ZDp������XZ��c���&�E��yɠ53%�յ�S}�7r�����0�>�Ia�Li8���l�a!aX����[YᏯ~&m͉��?�#�K�D~IcQ}E�Ѫ�4��1E�j��a�l�5�vG\�]��T��w�._�:Jw*ն-Z�7��.Z�N�e
Vl�j�j�U#:����b��,����r|���/&��+�&�d
����^T���w�X�#Ơͺ��ʵ�A����b�4!��Z\���qه�m�w���{��N'@����� �e�z�RP$I��
�n�ݡ�)�=m��t"ŏcְ��