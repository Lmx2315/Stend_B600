XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���#�w�9�ʞ�LY�W��i�����Af���^��������"�~3���s�eS	���ҙ�]���TaJ?�}�8D�$�G窫Q�g���Ū1��Rj`�[�~�.���)cZ[+��b6㋽�JQ�h;T(	a�d�Fc��wm���J���Qc/�[N �?�{Z�h�'�'�c��N��2�}�'2�yi�͂F��zzi������Mt�@���].��q�Hyq��3+F� �6j�`SA��n�Q�� W���*6tt���ڵ���^E���%��=GF�j�gl�<�J} SQ�n�R�^�Z�t�+2؏an��[��3o< ���)���9b%z{�'ncj�/�lK�m����iUg��Pk�c��􈈯��j`�gր �W|֛���(w�p�$��)�ᒍ��N%��uC;�j�|�XU���8jY�	���R���ԓ��[N��^���qt\����<� :GgI�,b�s�]�Vȕ��S�(���l�Qu��UP�����z��ge�ܮJ6�������ھ{�j=İ�Ьz�g�l؊��@ȇ«i�OƐ�j�k�#�ǩ7WFn봘���Q6{��1��'��슐�W �pT���wo�'O�uV/��lW6���v���"].���t��T��`�������@F�Q��|b��*������l>n�+��s]���	��6�r��y�[9ӌO!���7C�&��׋�+�_Փ��=<�ѭ��$�\�^#JǀK���3���XlxVHYEB    6fd8     c30��n`�ɧm�l�3dܪ�?����o���?�_��1+A螼g���6�ٽYAJ?LKF�;�#�DR"���KFUJ�^F ��J~|���nFf+�����.*�/���ǝJw�I�V�g�X��t��ڢ��zK��4��Po<`磨����$Â �G�g@�tT�4\k�=��!H<O�,x ��TF�6=f�su��!EƤ��*(�_�s���53;��c��-�@�s��d�)K�"��=�ՅN����	),�*��;���k=���u��+b��*�HG}���D`b�= ����*�]#W��	���c��0D�3G%N��\�V˧��`�����ߺVP��7ФO��껐�aF�mtJĺ�������~��ԧm��Ũ�_�v��z��i�FI����������b��a��p'�hF�pɈ x��p�()>
���BRRzJ�{U�g�!�T��|���#n�e��z����]��nk� ���xe��5���l���|c��ש=\�v�=�����	]�\���h_i,6�8��*|�ᨃ���=��0��e=͆Jt8�ݞ����� I�}���ö���1(�ըZ@���*��?�����{�$W\Q闛I�7�_05+c���a"DR�_�V"#5�v�5�2�i?�Ғ.
�P�Y�mY��NU��b۸�\�����Ru�wނ'҃�h�L{�+	�ؒ��m7�
^�Z@���(	�ü����([�w�}K��+Ŵ�.�/WU�M'j�������>|� ���d�R��9�/��XӚ�����F�Z���=m�9��g�A�h��K'���5�L5Q�t�Թó6�Գ���o�����M���nضg4��o]�T���ʭ�&Rf�k2����U~��X� 3q����=���KO8�]q��V����UO<�����V1�[�k��x�*,MM��LY�'�l��!��� E0����B�n��iv�V��
Rf��-��N}�bB 2.�D���A�ǌ'I�;�SE �%��ɖ�Ug|���3oNG�h%-K�Vl�ܮl+����YҢ�cu�D�y�[)��5��6{��"4��Yr�b������c�r���p;&i��;�6}�|�+�����{T�eG���v�{�N�ŵ������EӯxF7`�\��a�[0#*¦˘�.ku��x��V��%��CJ�5��Dk΄_�K:�Ӵ�����hd��T�2�*j#���7�vmE�M��I��n[�����hX;3ӱEs.O��Z����|����)L�=��޷pk�A�h�Z:�����뇉���8�{ؽ�v�rIFݟ6�o�l�jjH�v}-�<�=�y*B�&E7��\��������װ�@�1����I�R@_N�=�d�z6���W�U�������� �Q1�W{j��n�`\G�E���8�� �v�B���/- gbbt�)�>ԑ��Tm%������n�#vbI&�4=v�b�?����p����2�����dʜ�Ve�n���X������>��q_��(<_Ѕ��O�{�]���;�%��7�����~Dĝ#O�1��A$�xP������O����r:Ջ�Da��*օ�:��X���f�z	��/�8"��Lk��OT?*�k� �Uq���IN���?Ll�	rh�����x;��o�;���^���[|�4�5=3d`\<�ǥ (�lzK��C.�~������f�y���5Rg��l�'�Dn��u������5�d��R�!�?�(�NN����n�@>��H �s���1���ء�C��i9u1���"G�f��QA�ʜ�`,�q4�_/��H[�VD�v2סDH�9/j�YNM��	4�("�/�lB��ꌎkrɧZ�(���7���Ғ)�$��:�t�l�.�,�a�S�:Q$O���{�XB?�~�=6��*a��	 �����l7�������Ԍ�h�J�ۘ�)K@`�O����E�u�|�.BC�
G�U��i�H�	bH9{5��MHfM��G�z�����1���N�Oa��S~�*V?Sz�Ov��ت{4�Z���L<�����CZ5)~MP���Eh+#%dW�Ѹ@&mu{c˸����\@�Z[Z���k��'���I�3Kz^�*T|i;3�d`�;��`�Ӧ����;�Yq��i߶�׹���TkJ&�֎:Q�e�v�A)F���T���/1�k�lZ/S�qD��>N�� �:~2���Nc�~+��K�4�L�i A�S2��}�R��:>E��N&UhE�]q�����^�� k�G���}���B�֮����?<N̡N�Hl��-�QNR(l�vl���A�iB �4�(i���!+Br� E��hr��%���c%s����Ũݺ�ڶ���H6�h�%,l*F`��س�{�Q����b�n ;wOq��=bp�-3�8ТZ/l�{M&0h)��iNr\֗9k�a��X��W� �c䖐``���9YD��
�m��)���c���Q�r�g��aP�	�m=7�Tb�ߝ�2�-�x8���R-��.�HD���i��M�NM^��������:A��v
s�M�{�?<�����
,�)_�fJlǨ)Y���r�0������x�d�uQ�Q*�9ye�Ѻ��$ƃ��0���"��+<T�$ys%��+�.�S��2M�lV&_�E�B�'X/X4 ��l��t����aw#��p���3C��M���zp�-W�<�[���C9����>3g591�l�snk�&�n��J�"O�����M�pS~���;���BS�nplQ��Ai2%!kn���l+y%dc1-�A���Xq�Y���S�-.�i_|&5��~���Km&m�;p���_:��H�$$��6$��CI���-\T�G8BO��ڛ�#�=�+�Uj�Q���5�A�D��,}��K����h������K����6ؗ�F���U�IE�0`���~�0i��-��Bg�5k$��7���7�zvG��C���Z!q;L�t���3Ω�ٛ#WH.c~����N\�X�p�鱜�i�GTh�/��ag0~k�Gɳp��