XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���r�w�۔��p>��֝�'7e����5���-�7qu6���]�b���Ub0�S���	�<�Kz3UY�~�g�ڵ���n��r�Q&�`*�I۳L�����TS��������Q&��/��yMՀORy�l�"�,;3;�f���p�Ƚ��QP�5���6��'����U���TT)(G9��	>�������c>���&M����b��O�n
:��_�۔�V����rè�����}��WD
[xT������2�Jl2}�>�윙��N�#|X�W\I�q�����Ou�X�r1,�2�j��~\���=LqSU�⌎�dE��35�>��bXoQ(�Y>ď�c��$o��5R�%eX{���mVй�2�m����{�ꐀn���v:M{���l6�
�NdM��+���k�x~�ط4�K�����9�]�\�p�Ý��x"�_?�xOwʫ�!�������upG/-"�M�n���QO�Vah,ݍ���s�N��Do���h=��~�!<�Q7+��>�������lN$�p:d_c�d`����M.�H73�W�����\�-=o>�H���A��F�EyG31��i[}���V:�4�@��s�������FF�h5@��q#�;�1 !�C�=�	S��.�t��'ڔ �HT3�̇�	 �C+Ԯ����x=�61SGT��\Cm�"!Aӛ�[��;�х3jL��_���րl�Ml����)'�P��b���
J�>���e����7nS���O�e�+VXlxVHYEB    2d5f     800I	�#d���Tփ�*��ah��wG�A���N�:�6�$Oz�[g�8�����q�/�2<�4����[w{m1�4�~W�K�Ѻ��j��^�i�#w���G폔����)3��GŬ�������L�MA�8M���w�6�� �p'z_V@�aÚ<������в1dX�]�8�GH�*\�$6A��&�8�}h�FD[d}y���doZ �u���cլu�P��)�����j�S��*?��H�0���V��S�����Nv��+O@���6�Q�xJ�.��X�T������JK��̰�m2���z���yV��kē��	�T8�dd�;��+A����Q��*�*�� �W\\��E��"1���8�B�۾��O�,��lX&N�����|B?����=��w�-Rԍt�%?�L��Ƒ�I5�	�<vɒ�HY-9��Z8-˛��v�b�{_�@[���/[w�;J�펍,�� ?н�W!����� @gM�"�ڵj�R�Bu&���o�S=���7���xPC�2�Q%p��?�G��I3J9�E�l��&��3�y�K
����v��cbPhz��ft^T�u���@���&�ZR������w���V"�0�b���nx�sy&�Ch5)�� �����:��D�P�Ցm�,�e��W�;�?�G��Ȇ���Z�S�m�
҈����/nÞ����� �]`�B��y.&Jx�w�4GV��Q�J��o��2�o����O�-%bHJ� '2Km%1�̝�Z����-���?�>�����A�M��Y�ŭ�7Q�������Ȝ�d�1<y�$�n�`J�FK�M!�֖�:{�@�!���]È��9�2�9PZ��*��v����/&���s4�$# qz�}�S�--�U݇�;�԰4��.ϊ�ZGo��j-]z���k�Ɛ�*�W��8�٨�^P�D�2$��)��M`̹X������a��lH�
WA^۸��降k�1�ʔ��$B�{�"�9�Ck�F؎j��j���ސ'6Ph�&��G��΄:n������V�y����}���z�n����]�!�3�B8MpO��S&��q�ׇ��nw���������|4��2,� 띉�Gy�6KBڒp��ƽh�a*ĵe �X�T��<�� ^�A���1���)�>�b�W�ǐ��R N^!�4nV��W�������\��7�K�����_� �eb�@�;�ؾr�
Q�\��Y�>�r�v'��ΖX&��>��B�g&gb����a���/f�vȅ��r�Z�8Fw� �Ntg�x�~�swz�������{n�������_���!���$�4㝚�3��p��v��az:͇R��q�u0��"�e>/²��(��H��x�U�{p`����]ˡ��+��&%�'E�]����RA��jN����@D����6B�,��>�S�qS/�:;%�������㏹]�d�Rha܌����-7��k�<e�,���F,ֲ
b�Z�ƀ���7�j�Ġ�L���Np�J�\n(��!̇�Ϡ�g�3���؛mQ�(��Z,����a_E޾>&�-���j�Ҕ�c���U�6w�N����s�IvPf~���d60��f�Dw�f����?Ay���mx�g9��k 
��n�6yt"I�X���z6y+��'琕Zg6��½�7kԹq�&��a1o�7�\���?�GJ�6���=��B�T��U��Ep��L�;�t�0n�c�"5e���0R�z�����xJrӔ1����+`ӹ.G&A��/��c�"=����|};~�@9��G?�0j�bd������0�3Q�g�;w���6�8�������<�N�d8����B~g[zn�^��4R[�]g��]���};�X�JT:�^I����ί�?�V�ip��խ9��p\�4[�d#?�V��z��cj�=m�%,� ���t��zl|Cu�������C^w":@��t3���*&����	�1����
�U�X$�љjR[