XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���#3��q�F4�š�M�nbF?�Σ]므0J �e��Ql�H��J��bX#��Dz�<��Q��l������h9&y��V8+����r~Yb����aJ��}O�)g&K0�AO �|���cSF��0���Ұ}e^�֎h"Uv̀*yZ��	m�Hxo|�������Ǩ9���҂K���K��bpmӒ���	���@X, ��g�=E�('��e�Hq�B*��Mm/H�&*����L)-��A��H��G���X�ia�Y��4~q�5�\��FoQ�*;�N�\�S�&A�Y\]��
�9@�1��.��v���-���K����R8ބ��pM_H�n<n������w��B�izu�e���?B����?�Ֆ��S���y��W�%)��<�����i_P
ɒ�Q�B�ه�|A]�I����)�X5�sE�%#�H[!���.�t(ŏ��Ƙ$-��l��A�#���Emr?���B���AO	+�O�q��I��Mп��EM�u\��JZ���7���,N�MuE�ۨ���UF�4�B<F����J�v_�-�q0������"锨�h�Vv�n�r� c~(e�&ڼ�ַ�K;X4�����Y�}�L��^z�]�8B�oLʪ�?M]����@m�q~���@�NY�M��Xģb_KQ`��&����HL�Q��ҺyV��h��&Az�����
m}��?���d� �l�M|��Hi��1q�������S�%� 'Ղ���Q*�,K�߽ƽ�q0�ҍXlxVHYEB    225f     610O%L�F˘��W�軚B�Y91:	\u&(pٚ���(�I�1���Õ��QtXr>�W@^��a���X��tu<cceˬ7hta�3+���h�
�b�ַ'7�ڙ�џ�7ݡ!1�%�d�1F�-A�����d{�3�E�B�?�k�V�:��JWHn��$t-�$�ܙ��MNlȮx8�2f�&��g"M�$d��ɡ*��s�8�_*�I(�J([~{h������-u�TNM�ï_l��b7w���1Wl�f�Q۞���(�����h�:`��ex��<����	��p{�X�X��#C�����$�w�
rW+!9;vA�կm�t�!B�Lm��U��*&�w��F*��u� Y��ϣ&��r�G�!��Eyy��A�+a�Z�(�A��|��XY0J��[��p�n>�����4l�����Uf����ﵚ웵-`���`VtS��+�:��\1G�8{j7w! �p@`[5�bi��Z@����2f3مS�hj�c0��PVH�3�ǁ>Ear��'<"n��.e��6ߥߝ�y��jGX��H����N�B|�9�=�e8o���3�Q��e�4%����Z?X�lJ�e�}�m��g��%qLOe�r��Ĥ$�W�<c_���$���Ţ�0#tx�GL�;.�Tx��P�YN��=|]�f��aZ���Q��~�Q�A#w����em8�k��rt9[�I�I k�z�nϮ7w#�x�3@=$�x�4����Hd#ƊUCj��%�cݦ��j̠O����
�P-�N�z��4L�d�p��E���G��)(�yp��5�-]�`$h5�uK�kD�ŏ��)0 :��k��!�}0���+��`fb�τ�{�K��\��&#�r	uf���DX�qČ��a��:c�����A�0iF(j[���6��}"D�r̟�g��C��V�M�f��@�*�u8rgӿV��)��鴙�C�)y!�#ә�����t��ts��,<��py�ҒS�{;�?���,�/���� �����v ݖV����i��R0��x����N���v�m�ԎJ�z��p�AnmtӺ�K;ƨ�������M����?�Qݰ����`�����bf�Ub�����5כ|~�f�;��t[�N�ul�$]�
��ke��Jf�����}˫N���A�<��@���F$J��9�k���x|l��(�u������=�-�m�D�1{P�D?#
	=i�#4-#�ج�n"�r8��E��1����sc|0؎(�X���:ﲞ7�q�XF�o�:BS5�����-�2�.}�\%ݺ�pƮ �*Hr�Ɓq*J��_�>a2i�$�or=�k�p���6|P�2����D��YQ¾yM��ӾG���Fi���v�7�0{�Ů���.���Q�� F�7h77z[����˳�4�nK��`��+%8�{LG[�~L��n���C=��`��O�󔂖 �W_�{�9S�:[-<��e�/E�Lh'�ڡ������;�H��\�jV�'�pʯ��d��<Qb���]�{