XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��v��>��1JL�v��J����;r�P~1t�+�)g�0�
&�!���՚�[;�2��o1�I��b ~���1�X����ݣ�%u3���B[����ND��K�N���2�W����K����$������~=����!W��m�:��ßgծu�	BmzM��P�d����qC(T��c��O�vo�G�T&v��"�o�my�[��9�S�K`��y��π)���W�|��1Ί�;��I�u�_4v��eMu�_}�Z,�l#O:��4������Pؒ=ޠË��oM]�7iT�{�C�`�UTZCՃq��>�Gj;0w��գ�nE��o��/?ͪ��-�q�S�t��M�k[�*ː�a�ް,�Λ �x�9��u��%���{�ο.T��A{�p����+%����H��ޜ�v��qI��<����� ���}��84��$�DK���4�2c#3����:o��ƣ���� ���~��Y	�VVch��c��,Ak"m�k�`@�r4�}�q~lji�O�6[$X4�!������#``���a/�xB\j�pn�e	��P��Zddt���Fzi�G����2Pc}��8��ώc���j���Z�X���ZƥC��׭1f�ċz}�:�T1��  �tm�uQy����ٶ������pw?�8�5���\8K���Xj�	�5�Gz`�h�Odwv��ЭC��*�M��ʣ���h���r����K�%�j�=�]�g�1���d�Z�[XlxVHYEB    1577     5a0��@��@���ګ�9�o���^.p�8�+�0]|�V��s��(	w�>�����0�~��:�tWU!̂�cy�_�@ݜ��'���y o��1�a�����Х��>���K�A�Zk}c���<N*
�.έz1
?�j[f"����?8�l_��I?���X�"o��b���I=�4Q,���5an|���%,��0)^�C
?����Ad�2��.�eްGt䎐Y����cwdN��i�>y���ܲ����'#�D�����T� _������K�T7�!�x8��Y)���hK�"iD�z���r����湛e�(�ÙF��u��Q΁fc2�Gl��N�!S�*�X)w�H)�@�5��Oy9�FⵃBtou���y���3���*�G+�^xR�x4���	�O�9�MzN�Ϸr�ri�\����fځw{ j�f�	�X2hAC�P؞����<A�fؒ�i��<��˭�QУC��u�o,b	�)��Ö�����ٝ>�]j��f�?���@~�;i��m�G���A.����IG�rJ�^$��wW0�b�M�#�C-�tq�=�S<Y�ޖ�γ����%v�/�!���=i�v�X��<�m0ZYo�&��x�E�2!�q�d���H�R�$Es5����@K��l6]���n:_^�!7��y� ������l}�j�	*~U�L�$���S�KBў�@��Tr��������Qm}I^MCk�6p�N�e�O3������5s L:��WUa��vOER¹cWv=�vL�QC�t��T�X<�66�C	���3�In�?B��z�"L�iڲO�f^�xؙ��~W6�M9�v?׃��xd����pQ�ʬ4I61Ab���������B�w���G.a�K�fN_fs>\~����?�f�<���l���H` �W�`�̟�$��j��M�b���гOoُ�s���V�t���d23�7��f��z��$U�WMy��`��y*�d�v;E:\���? +�r��%�����(�ߵ�(���T�Z��Q�ͪ�,;;�B�m�.r���)w��������s�Ζ
���L��},,$�� 0?���a��*��e���kz�*8c<�;�e�3��H��"3�'��`�Â��g�g�i�hzc��eB�$57�m?;W؂o�X��V`"N�5�C�_p(��}H��3�e|z2�>��@��+zQZ�j�}mJ�����v�HQޜf{ f4��ї�IF;&q���Р7�aD9%���bs~��M��vc��K���x:��&;1����-����Bӹc���;�40��(�J�2jʈt{X�=T���/�y����G�����q��4͢�f Y�N"�c �Db���=2���^t���X zj