XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��3PTu{Ȏ����(�޹|t����g���}����X%.$s�Ƙ���$A˅��ix�BNyO��\lC��Zm������~@�;��k�̰s��&���=�}#jE�����q�lz�+W�׊ucD=��|6�Ѳx�=�'�~��旋����`,�A��Vr$	8�E��El��šO4[-�R�y��Đ�y���C�Q�*�s!��O��s��J�Z{��9��!p\$kFD��g��z�>�D��C�����)�4d�ȥPC �_�Bgy-��rF@�����N�0B&d���g���:�5|��q�o �|@��珬F���u��ŉ�����7�����#h��]�U�̸t*�gR���{,�����ʿٝ�k@Rf�z�s�r�t�T��Z�{v����[�c�mq	fq&m�P�_7"y��'�'K�o���Z����F_]͆�qU�+4-9���`9�ul�j^m�"�Sr�xv��s,q���!N��1�aZP4���zW�h���Q�
&����?OAƦ���:k�#�*y�J+�������,��D�!�/-��iJ�P��Ipۣ����e��R�|B��G3?NR[˭�Z�oS
��r���6ThI'6�$Ȳ�ׂv���8���,m	����[K�DY��h�[R��\�J ��{�� �������N�x�9��h<��Ť���Z$J�4��D��4�ꉫ�'��P +��-�&87�>@˽"%K��z�"\�e��Y0���˽ �XlxVHYEB    1047     4a0*V_
X�:���釿�ף�ěp)��|wDc�v���%�ګ��B���	3s��9'
}�i���_�ұ(Pl���WaI	��w��E��o`����mG�Yo�'sK����{
;E�w|��0���|�m�o5~�cY�N�翷��̢�֋�K��F8�O�`�.=����8|�	u%��9	6�C�s�>� �x,�����}�?�4���`�*f⪵A�O�<N0J8����Ϳ{����_Ɣ]�0�wX��	�K"���2�@^�*�Ou�%ɾ�n2�I�H��0�E2w!�1W��3޲Ӱ��r69�<����$��CEm�|h��A�f&��닸��RM��]�%�u:��[����=�Q�V}�<�Ȓ�/46�`�}���#>�y6~bʄr1q$�Zi՝�S���L�� ���BX�$|�J���H��@/����x~���*�F	��b���-��=���i_�����i�6�Q�~J3(E�y�G����P�Ҙ�T�B��e�y���f�V�Ri�y��C ]���"!7x���_y�j��۞�Y��X��
�[ǽw�Y����>�6�G�$ѾL.:!ҭ����yǃgR|y*��2�DQ�2�b$�S�sl����O����wpqj�(?sΦt:
z��i���([�V��1B��Pf<6%7�	i�	(����>�n��"6 �LTK�P����Z�3�O�hݒ��j��Ѕ{~��߿�5L[0�by o�Z�f*#o�줂sz_W�_�7�0G��K爏-{��ݞM�jx���б���;��6|��,��,��F��~����hl��_��$�=��)C{L����0�����F�l(����2z�bG`V�c�?X0n�e�KN!��ֵ��>�I2(t��SQR�ړ�̲�7U��wj��u��F��	D����{��,���w�?A�Qb�:e�O5�n�'�.���Ӵ��Ԩl.l5{����]N��G�d����Ӡl�Lc�8q=�2-Y�F�!W
����y:� |�gj/���#�~i���W\�-`���d�u���u��r���60���9n;Jۍ�4=��I:%�@�˃/RN�T��Ý�QyaK���]?A21E�D�㛮{���&[߳�b�Hj�d���]�3S�b��>��!D��